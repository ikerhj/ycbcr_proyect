��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.
zvߠM����l7_0� 6��<cH�
�'�3�H�������},}����U>�z-�?�\�7Q{��(�'�`����B��eHm�g�(`��v9���K�2V��*��("-�χ����,{���@LR�]���e�~���V��C�*�C;?��5�
���~,΃R�ssu�J$c�-uK*0��9��9�֒�e��%ߥ���l���8��>�m�^�q�x�"����1�u�|z!*�{=g�G�{�y���-�֭<��=�y��ށ�1��]gv�r1G����X0��`{�������71 Q!\'�/z�>����k`�%B+Q�s�)Ǟ�=H���2/�'�fd� ��h��T�Qn�d]^��ê���m�U�X#dI�nL}���� `��CM�Pg:��'!u&��"�v�2��[����[��N�$}�u�F:�Nɳ@i�pŜ��Ӑv>��S�ol�_�P`�ЫGxP��Î.�w0$�ɐc�t�7����:��e��aŮ�1)a�F)�(��IE�k�ͦ�(hn�3��j�n�����Ra�T��p<tLw  7�j�ܧ"s��'f�V8HL�Y�H<'6��hy����t*�\�|a�4�)��0�Epjo��waلxʒ�T�5G���~�:v�̦�,�n ��91��ɛ+yc͏�1[D��O��T�ttd�	p�P�IF^LL@��,���D��y�A��6KQ��&�ՈD#�E�A�啖��O]a,J��Gs�\�G������g�0��hO��Vʟ�3�%Ք
E(1
��!�4,&�6�D�&�����h̀�*���EZ탶�b5�����ᱣ��r�r�e���
l��2pB��>[�VE����V��ӄT�M���FS�5�,�ۋ�������>�+�œ�/x�eE-[��rA�*�ͫ�v*��9�����|��fE�<
#!�]�"x˦t����w�7z�	<�7lsl;��`<S�I�!��~+�[�ץ���t��q����l������wYȬ��d�i���]�A��܄<�t8�jo<|��	D�=j�л����S�#�gs�dM�C�������x����]i�,��hp�~%2�4�h@Zr�Ȁ
��@ �R8�����HX䠈xM �-5h�B����^G�hp���g6�A.��c�&�I��t?�Y��ăHX�D��0d�.�W���K�����_�M|�L	u��Q>�3���\9�v�٣�J�T�*��/��r��[܋�X*#�5&��t�_�r�ߑrO��b��op�d�q��>ne誈�^ݹLR��>�ϓ�k2K��PA�I@qM�/j����oߔp��Ud`踦�[e���+z����'�Y5��el���嶵Y���ꘂ�&W�a��͕'�^5`��Eok�F�Vp��F��0��s��aw��4��9�lX�Q0��vW3 ��s��E%��4�X]���t�ڷ!���m�璩&m�������Z>�򁜶S�B d �ئ%��'�`Z;�u����kY(�?��Q?��s�����J�J���K��6e�J��I��$�5�n�L>;�p���2��M#�	oh�T� 8(�Ŕ+\Bā�_ZǞ�Ml� ��C����!i,���;����S��x��gv�%+���*��O����P�/���y��w���%f!xp. �a�6߶���N�����Ui�G p;R:bM�]t�$̂?�N�����d��B�"� �F�"bE?{o�}ID������?�A�G��"������Ug�I#?��U�{$q%m��z�^	��������R��M�	�4��!ׇ�G��0�a�?-9�Y����e�M��<���#���TE��n�K���X�#"T�$d3��v*����ovv���e
�gO<��d��ꕥ�����̨��[��F+B�d�>��F���+�Κ�oNZ�������D��➢�GR)��U�E܁No9�a�3?�~
���=�[�'����9t���m�4�['�1�����[kN'ȤY��,����ER]*K	���ZU�������
��/�����.�+{�i��VM1� 0F{��t~��NH�e�g��������U/��k��ǔq8"�\�M�h��Y�_f V>Iq����SW0��?)��j�:���ثҔ\�	��y�YE�o}!�-*>Pk��wH���i�혵Ѫ�d��,�'�UI��K\���*ʽ�3#RA9�Q7�T{&&��]��>�F��lT��'�7��l�������ݞ1-s�Ep����h@�t�.���[Ğ��1���1�Bq_C&S�Сx�����a��K�T�s"���t9�D��E��%{S�L��>_�y�<�ꩁ�bk����9���ѫTrJ�:����JN���e�b�O�UZ�F
ǽ�.��px���*/)�w��
�'/��4�U�Z����d�qv$�T����CE�:�N�(��aձ�{��̵�Ώ��x5�
�2�y�$�jc�p�֊(�ׁF�'���'�5���1���]�{ CҠ�m�t��]��A�t���;�ABEwF�S~`$�Ѝ[�������I~P���}rw�Jn�3
ڇ������J����r��56��������	�?�x�ej@f�d6n0��RT%[w��շ5\��,Bx�K=A>���t��j鱭��}�sU�}j��|L�`�k��y�6�(����!�{4�8���P�Nd��<Ǚ�e8�>;/��j���ȽX�N"$�S�v S������y����-�Ը�\[<�ۃ�0�}$�Ok��E�,]1#��_R��,\k;�y[W#\�/�=&��U��q����<�F����a��'V�&�2��@s���M4.�:�8b>�1�R���D"��?��.H+���&����&oMl +�C�$�������4����}��������'i�۰C=��D��
QG^���]��nf����|*��/���G���lpA'�b4%�*͒1��P���ϭUw����{�C�>�ؼ#��^��2��ƚZ���t�����=Z�<;�T^<ZYIa�2��.h�J ����&�,�v#�_f7���p���q���_�t=r2+�Uj�x	�%8�g��� ��Qt.�#�'��9�Gw(�ƒ� ����P�MĄ���x0�u0:<��rՊ��ы����>o��ؾD���X������q/�a웯k�%G���p�d�ґM	�E��_��3!W�>˟Z�Fs���{����)�QpW,+�D���<�F���&=��}���7�C8>}92Q$ ��T��\N�Rf��_+�f;�1II�$y{�R#|�Ϟ�%Y�*���G-�*�c�i~�Y���9�P!o��߮��׺�x�ծ��/�������EW���"��J�r�@a�u�$2�&��+;�_� @��6���R�Q�0�}h �j7��գ4���1���4���>�E���	��=����qPG��,@���N�T��e�Dݣ9�Z���w$� ����!Я]�LL� �rf��翂ŕr�|l�x��/�
.O���j��H8+�&�͜�wW��Msˑ&Y;�����Ӽ� M�C�N)V�������AIFN�x��	I�B^�&D��u���C�뾇��ķ����!�r,&���<&H=��?!������;r���|�x��V�sR$�at�5�D��N2�"�C�X�@�7X�ƳP����@�b�/e�o�,y���O'����*%m�L����N��?@5�X���-
`ib�C��X�F����I�y���6�{$�g �Q���cs�hZ�!��j�6$|[�oG1�R�eIf�3񎮘������ߟ�"���^���������b���4U��fxn��d㯕�Q�R �ۄ��z[���PF8̤$i��<3W|%���*�d/���C�����!�/��G� �
\,�jN������9����hV�͟6�j��<7QO�|\��0����Aɏ"r�}[�v6�]�˕���[U����Z�j���>4K��2��o �|���4�w����K5�ڲ� ���U�����U�X���sNȮ9�<r#�8S�bg]�<�(3f��{z|E��`#F�LV*3���E�����K����a}vW/�:�5��g����Aa� C�a&�s�c����26||v�Ksw�����`-�NΡ	Xh��Χ��3����\ť~E��Ԟ��0cTfx�_>�kOA9����/A������Q�	�+K h�d�~1�jECX���^�#�튩�_���k��L5G�mo�V�C��9� d�T]�_�������J��W�~��p^�s�Ce��:��@§�XZ�K�S�5F)�&W�P��n�m��mO�7�����p{�$��88H�s�@	!݁p�'�q�)�5�f�ңLj�@�h����3O�M���f������AE<��_hv�c��E.�/���}�B0�?��r�t�QC��y������p��C��@�x�D�d'�1�bF�
Vj���&��/��^��YGXk�����p�1Q�a9=8��w��82�l������x(>��{�=��zI�v���_&!�������o�\���+,8��b��v�Ә}�������\m��u��a�:�w{H62�:~�) �r�U�>s7�8�C֧I��b�#?�3c}h�^���.b��ڏ�٠��a��E�#+y�	�r_�B�n�Ҵw*4�[��|Z���4A�bX�}�:c==�ڏZ�O��K?ց���Ä9�t�������g�xB{MĢ��ш�*��9�,�ӛ{�z>:��4uF�X���t�n5T���KMzuMNՉY�"�T�U�Wal�T�K�q����̮�/"������>��i��e�=ܜ�8�����2�h�^�Ù0Q�h~^M�����~�OeR�\[���]��5`>�Yչ�BwБ�*z��D����l\�o��6�Fk.w2W	��_�I� �1S�dILR�9�Ff�k�����G���t�xXT�x�k�]a�nՆ� 4�%���U��$JQ��_��A�7	�{�@X��Rii�3��~x���h����s�9o�妕�3�l�H��MC�?�#/�tX�����7�AI!=f�j�U�*)�+���-��;�����s��Nс1�u���j����FN}Ǹ�~}�.���!B]��P�B�yJk����>�1�1 ]H �,���H�x�l�x3kY�@���/�1w@�J��D�&N�zU|��eÔ���^[��%B�0����s��pQ�!O����ѡ6o�� �~��v
P9���K���p�.ß�q� PX�e}�h�D.l�f�SmRY�x��;f���(��usH�!"�S���0!�%�Ajxa���^��i^��BI�X�<��$3r��O��@�1�J�&�p	q���y�$�"xR��-�����07�0DG�X�v�oF/@��f8?wĔ�m��dN<(���ެ2�N���o�fV�p���屡r�E\զ�^�-�6��%���1�;Fy���� ��ep`��٬����DP�c5��럞��\�R8��$C��aK˵;Q0��y��$�J�촽5|g:���h\I��*�P��M��29������<�b�,�?|��̗'�zVw���\Rk%]Hws�/��t ��S�b��ƙ�X
�<��D]�^+s5/w-�_���g�����Tj�ei�A/E�$�f�RZgU�i�1�VC��YC����������2w�	u�.��.��q~�j]�B/��5���)C��![2㊣o,7�sh��X�O���>��h�G|�-?�jT<*�P)�X�O�����Ķ�0�؁vu����?�w�m��� N��Jlj=;5,�Y���6��).�WY�ɚt�ڈL?�M�a�̄�Ë�G�Ĺl���h%�nm��Hgh���Z̛�����T��� v�usT^a����sm��p1,,�^fh�x�wWDI�>���� �D������e袻]ľb���N\{@-3D>"�Xx�1m�2� G�E �<�S�BpI�X�^�$��>`K�A<nA��K���e������|�����
f�������sox��-ۓE�