// c5g_housekeeping.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module c5g_housekeeping (
		output wire        camera_pwdn_n_export,           //           camera_pwdn_n.export
		input  wire        clk_clk,                        //                     clk.clk
		input  wire        cpu_sync_in_export,             //             cpu_sync_in.export
		input  wire [15:0] hw_info_in_export,              //              hw_info_in.export
		output wire [1:0]  i2c_device_select_export,       //       i2c_device_select.export
		input  wire        i2c_master_scl_pad_i_export,    //    i2c_master_scl_pad_i.export
		output wire        i2c_master_scl_pad_o_export,    //    i2c_master_scl_pad_o.export
		output wire        i2c_master_scl_padoen_export,   //   i2c_master_scl_padoen.export
		input  wire        i2c_master_sda_pad_i_export,    //    i2c_master_sda_pad_i.export
		output wire        i2c_master_sda_pad_o_export,    //    i2c_master_sda_pad_o.export
		output wire        i2c_master_sda_padoen_o_export, // i2c_master_sda_padoen_o.export
		input  wire        interrupts_n_export,            //            interrupts_n.export
		output wire        mipi_reset_n_export,            //            mipi_reset_n.export
		input  wire        n_use_rgb2ycbcr_in_export,      //      n_use_rgb2ycbcr_in.export
		input  wire        pll_lock_states_export,         //         pll_lock_states.export
		input  wire        rst_reset_n                     //                     rst.reset_n
	);

	wire         nios2_gen2_0_custom_instruction_master_readra;                                  // nios2_gen2_0:D_ci_readra -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios2_gen2_0_custom_instruction_master_a;                                       // nios2_gen2_0:D_ci_a -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_gen2_0_custom_instruction_master_b;                                       // nios2_gen2_0:D_ci_b -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_gen2_0_custom_instruction_master_c;                                       // nios2_gen2_0:D_ci_c -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_c
	wire         nios2_gen2_0_custom_instruction_master_readrb;                                  // nios2_gen2_0:D_ci_readrb -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios2_gen2_0_custom_instruction_master_ipending;                                // nios2_gen2_0:W_ci_ipending -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_ipending
	wire   [7:0] nios2_gen2_0_custom_instruction_master_n;                                       // nios2_gen2_0:D_ci_n -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios2_gen2_0_custom_instruction_master_result;                                  // nios2_gen2_0_custom_instruction_master_translator:ci_slave_result -> nios2_gen2_0:E_ci_result
	wire         nios2_gen2_0_custom_instruction_master_estatus;                                 // nios2_gen2_0:W_ci_estatus -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_estatus
	wire  [31:0] nios2_gen2_0_custom_instruction_master_datab;                                   // nios2_gen2_0:E_ci_datab -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_dataa;                                   // nios2_gen2_0:E_ci_dataa -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_gen2_0_custom_instruction_master_writerc;                                 // nios2_gen2_0:D_ci_writerc -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_result;        // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_result
	wire         nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readra;        // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_readra -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_a;             // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_a -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_b;             // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_b -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readrb;        // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_c;             // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_c -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_estatus;       // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_ipending;      // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_datab;         // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_datab -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_dataa;         // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_writerc;       // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_n;             // nios2_gen2_0_custom_instruction_master_translator:comb_ci_master_n -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_result;         // nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readra;         // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_a;              // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_b;              // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readrb;         // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_c;              // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_estatus;        // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_ipending;       // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_datab;          // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_dataa;          // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_writerc;        // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_n;              // nios2_gen2_0_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_result; // nios_custom_instr_bitswap_0:result -> nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_datab;  // nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_bitswap_0:datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa;  // nios2_gen2_0_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_bitswap_0:dataa
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                              // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                           // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                           // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [17:0] nios2_gen2_0_data_master_address;                                               // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                            // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                                  // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                                 // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                             // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                                       // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                                    // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [17:0] nios2_gen2_0_instruction_master_address;                                        // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                           // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                       // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                    // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_i2c_master_avalon_slave_0_chipselect;                         // mm_interconnect_0:i2c_master_avalon_slave_0_chipselect -> i2c_master:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_master_avalon_slave_0_readdata;                           // i2c_master:wb_dat_o -> mm_interconnect_0:i2c_master_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_master_avalon_slave_0_waitrequest;                        // i2c_master:wb_ack_o -> mm_interconnect_0:i2c_master_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_master_avalon_slave_0_address;                            // mm_interconnect_0:i2c_master_avalon_slave_0_address -> i2c_master:wb_adr_i
	wire         mm_interconnect_0_i2c_master_avalon_slave_0_write;                              // mm_interconnect_0:i2c_master_avalon_slave_0_write -> i2c_master:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_master_avalon_slave_0_writedata;                          // mm_interconnect_0:i2c_master_avalon_slave_0_writedata -> i2c_master:wb_dat_i
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                        // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;                     // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;                     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;                      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                               // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                 // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                  // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                               // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                    // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                    // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_hw_info_in_s1_readdata;                                       // hw_info_in:readdata -> mm_interconnect_0:hw_info_in_s1_readdata
	wire   [1:0] mm_interconnect_0_hw_info_in_s1_address;                                        // mm_interconnect_0:hw_info_in_s1_address -> hw_info_in:address
	wire  [31:0] mm_interconnect_0_ext_int_n_s1_readdata;                                        // ext_int_n:readdata -> mm_interconnect_0:ext_int_n_s1_readdata
	wire   [1:0] mm_interconnect_0_ext_int_n_s1_address;                                         // mm_interconnect_0:ext_int_n_s1_address -> ext_int_n:address
	wire  [31:0] mm_interconnect_0_cpu_sync_in_s1_readdata;                                      // cpu_sync_in:readdata -> mm_interconnect_0:cpu_sync_in_s1_readdata
	wire   [1:0] mm_interconnect_0_cpu_sync_in_s1_address;                                       // mm_interconnect_0:cpu_sync_in_s1_address -> cpu_sync_in:address
	wire         mm_interconnect_0_i2c_device_select_s1_chipselect;                              // mm_interconnect_0:i2c_device_select_s1_chipselect -> i2c_device_select:chipselect
	wire  [31:0] mm_interconnect_0_i2c_device_select_s1_readdata;                                // i2c_device_select:readdata -> mm_interconnect_0:i2c_device_select_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_device_select_s1_address;                                 // mm_interconnect_0:i2c_device_select_s1_address -> i2c_device_select:address
	wire         mm_interconnect_0_i2c_device_select_s1_write;                                   // mm_interconnect_0:i2c_device_select_s1_write -> i2c_device_select:write_n
	wire  [31:0] mm_interconnect_0_i2c_device_select_s1_writedata;                               // mm_interconnect_0:i2c_device_select_s1_writedata -> i2c_device_select:writedata
	wire         mm_interconnect_0_camera_pwdn_n_s1_chipselect;                                  // mm_interconnect_0:camera_pwdn_n_s1_chipselect -> camera_pwdn_n:chipselect
	wire  [31:0] mm_interconnect_0_camera_pwdn_n_s1_readdata;                                    // camera_pwdn_n:readdata -> mm_interconnect_0:camera_pwdn_n_s1_readdata
	wire   [1:0] mm_interconnect_0_camera_pwdn_n_s1_address;                                     // mm_interconnect_0:camera_pwdn_n_s1_address -> camera_pwdn_n:address
	wire         mm_interconnect_0_camera_pwdn_n_s1_write;                                       // mm_interconnect_0:camera_pwdn_n_s1_write -> camera_pwdn_n:write_n
	wire  [31:0] mm_interconnect_0_camera_pwdn_n_s1_writedata;                                   // mm_interconnect_0:camera_pwdn_n_s1_writedata -> camera_pwdn_n:writedata
	wire         mm_interconnect_0_mipi_reset_n_s1_chipselect;                                   // mm_interconnect_0:mipi_reset_n_s1_chipselect -> mipi_reset_n:chipselect
	wire  [31:0] mm_interconnect_0_mipi_reset_n_s1_readdata;                                     // mipi_reset_n:readdata -> mm_interconnect_0:mipi_reset_n_s1_readdata
	wire   [1:0] mm_interconnect_0_mipi_reset_n_s1_address;                                      // mm_interconnect_0:mipi_reset_n_s1_address -> mipi_reset_n:address
	wire         mm_interconnect_0_mipi_reset_n_s1_write;                                        // mm_interconnect_0:mipi_reset_n_s1_write -> mipi_reset_n:write_n
	wire  [31:0] mm_interconnect_0_mipi_reset_n_s1_writedata;                                    // mm_interconnect_0:mipi_reset_n_s1_writedata -> mipi_reset_n:writedata
	wire  [31:0] mm_interconnect_0_pll_lock_states_s1_readdata;                                  // pll_lock_states:readdata -> mm_interconnect_0:pll_lock_states_s1_readdata
	wire   [1:0] mm_interconnect_0_pll_lock_states_s1_address;                                   // mm_interconnect_0:pll_lock_states_s1_address -> pll_lock_states:address
	wire  [31:0] mm_interconnect_0_n_use_rgb2ycbcr_s1_readdata;                                  // n_use_rgb2ycbcr:readdata -> mm_interconnect_0:n_use_rgb2ycbcr_s1_readdata
	wire   [1:0] mm_interconnect_0_n_use_rgb2ycbcr_s1_address;                                   // mm_interconnect_0:n_use_rgb2ycbcr_s1_address -> n_use_rgb2ycbcr:address
	wire         irq_mapper_receiver0_irq;                                                       // i2c_master:wb_inta_o -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                       // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                           // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                                 // rst_controller:reset_out -> [camera_pwdn_n:reset_n, cpu_sync_in:reset_n, ext_int_n:reset_n, hw_info_in:reset_n, i2c_device_select:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mipi_reset_n:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, n_use_rgb2ycbcr:reset_n, nios2_gen2_0:reset_n, onchip_memory2_0:reset, pll_lock_states:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                             // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                                         // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                             // rst_controller_001:reset_out -> [i2c_master:wb_rst_i, mm_interconnect_0:i2c_master_clock_reset_reset_bridge_in_reset_reset]

	c5g_housekeeping_camera_pwdn_n camera_pwdn_n (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_camera_pwdn_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_camera_pwdn_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_camera_pwdn_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_camera_pwdn_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_camera_pwdn_n_s1_readdata),   //                    .readdata
		.out_port   (camera_pwdn_n_export)                           // external_connection.export
	);

	c5g_housekeeping_cpu_sync_in cpu_sync_in (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_cpu_sync_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_cpu_sync_in_s1_readdata), //                    .readdata
		.in_port  (cpu_sync_in_export)                         // external_connection.export
	);

	c5g_housekeeping_cpu_sync_in ext_int_n (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_ext_int_n_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ext_int_n_s1_readdata), //                    .readdata
		.in_port  (interrupts_n_export)                      // external_connection.export
	);

	c5g_housekeeping_hw_info_in hw_info_in (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_hw_info_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_hw_info_in_s1_readdata), //                    .readdata
		.in_port  (hw_info_in_export)                         // external_connection.export
	);

	c5g_housekeeping_i2c_device_select i2c_device_select (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_i2c_device_select_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_device_select_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_device_select_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_device_select_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_device_select_s1_readdata),   //                    .readdata
		.out_port   (i2c_device_select_export)                           // external_connection.export
	);

	i2c_opencores i2c_master (
		.wb_clk_i     (clk_clk),                                                 //            clock.clk
		.wb_rst_i     (rst_controller_001_reset_out_reset),                      //      clock_reset.reset
		.wb_adr_i     (mm_interconnect_0_i2c_master_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i     (mm_interconnect_0_i2c_master_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o     (mm_interconnect_0_i2c_master_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i      (mm_interconnect_0_i2c_master_avalon_slave_0_write),       //                 .write
		.wb_stb_i     (mm_interconnect_0_i2c_master_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o     (mm_interconnect_0_i2c_master_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o    (irq_mapper_receiver0_irq),                                // interrupt_sender.irq
		.scl_pad_i    (i2c_master_scl_pad_i_export),                             //        scl_pad_i.export
		.scl_pad_o    (i2c_master_scl_pad_o_export),                             //        scl_pad_o.export
		.scl_padoen_o (i2c_master_scl_padoen_export),                            //       scl_padoen.export
		.sda_pad_i    (i2c_master_sda_pad_i_export),                             //        sda_pad_i.export
		.sda_pad_o    (i2c_master_sda_pad_o_export),                             //        sda_pad_o.export
		.sda_padoen_o (i2c_master_sda_padoen_o_export)                           //     sda_padoen_o.export
	);

	c5g_housekeeping_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	c5g_housekeeping_camera_pwdn_n mipi_reset_n (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_mipi_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mipi_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mipi_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mipi_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mipi_reset_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_reset_n_export)                           // external_connection.export
	);

	c5g_housekeeping_cpu_sync_in n_use_rgb2ycbcr (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_n_use_rgb2ycbcr_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_n_use_rgb2ycbcr_s1_readdata), //                    .readdata
		.in_port  (n_use_rgb2ycbcr_in_export)                      // external_connection.export
	);

	c5g_housekeeping_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_result                         (nios2_gen2_0_custom_instruction_master_result),              // custom_instruction_master.result
		.D_ci_a                              (nios2_gen2_0_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (nios2_gen2_0_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (nios2_gen2_0_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (nios2_gen2_0_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (nios2_gen2_0_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (nios2_gen2_0_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (nios2_gen2_0_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (nios2_gen2_0_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (nios2_gen2_0_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (),                                                           //                          .clk
		.E_ci_multi_reset                    (),                                                           //                          .reset
		.E_ci_multi_reset_req                (),                                                           //                          .reset_req
		.W_ci_estatus                        (nios2_gen2_0_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (nios2_gen2_0_custom_instruction_master_ipending)             //                          .ipending
	);

	bitswap_qsys nios_custom_instr_bitswap_0 (
		.dataa  (nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // s1.dataa
		.datab  (nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //   .datab
		.result (nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_result)  //   .result
	);

	c5g_housekeeping_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	c5g_housekeeping_cpu_sync_in pll_lock_states (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_pll_lock_states_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pll_lock_states_s1_readdata), //                    .readdata
		.in_port  (pll_lock_states_export)                         // external_connection.export
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_gen2_0_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_gen2_0_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (nios2_gen2_0_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (nios2_gen2_0_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (nios2_gen2_0_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (nios2_gen2_0_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (nios2_gen2_0_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (nios2_gen2_0_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (nios2_gen2_0_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (nios2_gen2_0_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (nios2_gen2_0_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (nios2_gen2_0_custom_instruction_master_ipending),                           //               .ipending
		.ci_slave_estatus          (nios2_gen2_0_custom_instruction_master_estatus),                            //               .estatus
		.comb_ci_master_dataa      (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_done       (),                                                                          //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                      //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                      //    (terminated)
		.ci_slave_multi_result     (),                                                                          //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                               //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                                  //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                                  //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                                  //    (terminated)
		.multi_ci_master_clk       (),                                                                          //    (terminated)
		.multi_ci_master_reset     (),                                                                          //    (terminated)
		.multi_ci_master_clken     (),                                                                          //    (terminated)
		.multi_ci_master_reset_req (),                                                                          //    (terminated)
		.multi_ci_master_start     (),                                                                          //    (terminated)
		.multi_ci_master_done      (1'b0),                                                                      //    (terminated)
		.multi_ci_master_dataa     (),                                                                          //    (terminated)
		.multi_ci_master_datab     (),                                                                          //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                                      //    (terminated)
		.multi_ci_master_n         (),                                                                          //    (terminated)
		.multi_ci_master_readra    (),                                                                          //    (terminated)
		.multi_ci_master_readrb    (),                                                                          //    (terminated)
		.multi_ci_master_writerc   (),                                                                          //    (terminated)
		.multi_ci_master_a         (),                                                                          //    (terminated)
		.multi_ci_master_b         (),                                                                          //    (terminated)
		.multi_ci_master_c         ()                                                                           //    (terminated)
	);

	c5g_housekeeping_nios2_gen2_0_custom_instruction_master_comb_xconnect nios2_gen2_0_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_gen2_0_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (1)
	) nios2_gen2_0_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_gen2_0_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_gen2_0_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (),                                                                               // (terminated)
		.ci_master_readra    (),                                                                               // (terminated)
		.ci_master_readrb    (),                                                                               // (terminated)
		.ci_master_writerc   (),                                                                               // (terminated)
		.ci_master_a         (),                                                                               // (terminated)
		.ci_master_b         (),                                                                               // (terminated)
		.ci_master_c         (),                                                                               // (terminated)
		.ci_master_ipending  (),                                                                               // (terminated)
		.ci_master_estatus   (),                                                                               // (terminated)
		.ci_master_clk       (),                                                                               // (terminated)
		.ci_master_clken     (),                                                                               // (terminated)
		.ci_master_reset_req (),                                                                               // (terminated)
		.ci_master_reset     (),                                                                               // (terminated)
		.ci_master_start     (),                                                                               // (terminated)
		.ci_master_done      (1'b0),                                                                           // (terminated)
		.ci_slave_clk        (1'b0),                                                                           // (terminated)
		.ci_slave_clken      (1'b0),                                                                           // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                           // (terminated)
		.ci_slave_reset      (1'b0),                                                                           // (terminated)
		.ci_slave_start      (1'b0),                                                                           // (terminated)
		.ci_slave_done       ()                                                                                // (terminated)
	);

	c5g_housekeeping_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                      (clk_clk),                                                     //                                    clk_0_clk.clk
		.i2c_master_clock_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // i2c_master_clock_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                              //     nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                   (nios2_gen2_0_data_master_address),                            //                     nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest               (nios2_gen2_0_data_master_waitrequest),                        //                                             .waitrequest
		.nios2_gen2_0_data_master_byteenable                (nios2_gen2_0_data_master_byteenable),                         //                                             .byteenable
		.nios2_gen2_0_data_master_read                      (nios2_gen2_0_data_master_read),                               //                                             .read
		.nios2_gen2_0_data_master_readdata                  (nios2_gen2_0_data_master_readdata),                           //                                             .readdata
		.nios2_gen2_0_data_master_write                     (nios2_gen2_0_data_master_write),                              //                                             .write
		.nios2_gen2_0_data_master_writedata                 (nios2_gen2_0_data_master_writedata),                          //                                             .writedata
		.nios2_gen2_0_data_master_debugaccess               (nios2_gen2_0_data_master_debugaccess),                        //                                             .debugaccess
		.nios2_gen2_0_instruction_master_address            (nios2_gen2_0_instruction_master_address),                     //              nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest        (nios2_gen2_0_instruction_master_waitrequest),                 //                                             .waitrequest
		.nios2_gen2_0_instruction_master_read               (nios2_gen2_0_instruction_master_read),                        //                                             .read
		.nios2_gen2_0_instruction_master_readdata           (nios2_gen2_0_instruction_master_readdata),                    //                                             .readdata
		.camera_pwdn_n_s1_address                           (mm_interconnect_0_camera_pwdn_n_s1_address),                  //                             camera_pwdn_n_s1.address
		.camera_pwdn_n_s1_write                             (mm_interconnect_0_camera_pwdn_n_s1_write),                    //                                             .write
		.camera_pwdn_n_s1_readdata                          (mm_interconnect_0_camera_pwdn_n_s1_readdata),                 //                                             .readdata
		.camera_pwdn_n_s1_writedata                         (mm_interconnect_0_camera_pwdn_n_s1_writedata),                //                                             .writedata
		.camera_pwdn_n_s1_chipselect                        (mm_interconnect_0_camera_pwdn_n_s1_chipselect),               //                                             .chipselect
		.cpu_sync_in_s1_address                             (mm_interconnect_0_cpu_sync_in_s1_address),                    //                               cpu_sync_in_s1.address
		.cpu_sync_in_s1_readdata                            (mm_interconnect_0_cpu_sync_in_s1_readdata),                   //                                             .readdata
		.ext_int_n_s1_address                               (mm_interconnect_0_ext_int_n_s1_address),                      //                                 ext_int_n_s1.address
		.ext_int_n_s1_readdata                              (mm_interconnect_0_ext_int_n_s1_readdata),                     //                                             .readdata
		.hw_info_in_s1_address                              (mm_interconnect_0_hw_info_in_s1_address),                     //                                hw_info_in_s1.address
		.hw_info_in_s1_readdata                             (mm_interconnect_0_hw_info_in_s1_readdata),                    //                                             .readdata
		.i2c_device_select_s1_address                       (mm_interconnect_0_i2c_device_select_s1_address),              //                         i2c_device_select_s1.address
		.i2c_device_select_s1_write                         (mm_interconnect_0_i2c_device_select_s1_write),                //                                             .write
		.i2c_device_select_s1_readdata                      (mm_interconnect_0_i2c_device_select_s1_readdata),             //                                             .readdata
		.i2c_device_select_s1_writedata                     (mm_interconnect_0_i2c_device_select_s1_writedata),            //                                             .writedata
		.i2c_device_select_s1_chipselect                    (mm_interconnect_0_i2c_device_select_s1_chipselect),           //                                             .chipselect
		.i2c_master_avalon_slave_0_address                  (mm_interconnect_0_i2c_master_avalon_slave_0_address),         //                    i2c_master_avalon_slave_0.address
		.i2c_master_avalon_slave_0_write                    (mm_interconnect_0_i2c_master_avalon_slave_0_write),           //                                             .write
		.i2c_master_avalon_slave_0_readdata                 (mm_interconnect_0_i2c_master_avalon_slave_0_readdata),        //                                             .readdata
		.i2c_master_avalon_slave_0_writedata                (mm_interconnect_0_i2c_master_avalon_slave_0_writedata),       //                                             .writedata
		.i2c_master_avalon_slave_0_waitrequest              (~mm_interconnect_0_i2c_master_avalon_slave_0_waitrequest),    //                                             .waitrequest
		.i2c_master_avalon_slave_0_chipselect               (mm_interconnect_0_i2c_master_avalon_slave_0_chipselect),      //                                             .chipselect
		.jtag_uart_0_avalon_jtag_slave_address              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                             .write
		.jtag_uart_0_avalon_jtag_slave_read                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                             .read
		.jtag_uart_0_avalon_jtag_slave_readdata             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                             .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                             .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                             .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                             .chipselect
		.mipi_reset_n_s1_address                            (mm_interconnect_0_mipi_reset_n_s1_address),                   //                              mipi_reset_n_s1.address
		.mipi_reset_n_s1_write                              (mm_interconnect_0_mipi_reset_n_s1_write),                     //                                             .write
		.mipi_reset_n_s1_readdata                           (mm_interconnect_0_mipi_reset_n_s1_readdata),                  //                                             .readdata
		.mipi_reset_n_s1_writedata                          (mm_interconnect_0_mipi_reset_n_s1_writedata),                 //                                             .writedata
		.mipi_reset_n_s1_chipselect                         (mm_interconnect_0_mipi_reset_n_s1_chipselect),                //                                             .chipselect
		.n_use_rgb2ycbcr_s1_address                         (mm_interconnect_0_n_use_rgb2ycbcr_s1_address),                //                           n_use_rgb2ycbcr_s1.address
		.n_use_rgb2ycbcr_s1_readdata                        (mm_interconnect_0_n_use_rgb2ycbcr_s1_readdata),               //                                             .readdata
		.nios2_gen2_0_debug_mem_slave_address               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //                 nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                             .write
		.nios2_gen2_0_debug_mem_slave_read                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                             .read
		.nios2_gen2_0_debug_mem_slave_readdata              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                             .readdata
		.nios2_gen2_0_debug_mem_slave_writedata             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                             .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                             .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                             .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                             .debugaccess
		.onchip_memory2_0_s1_address                        (mm_interconnect_0_onchip_memory2_0_s1_address),               //                          onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                          (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                             .write
		.onchip_memory2_0_s1_readdata                       (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                             .readdata
		.onchip_memory2_0_s1_writedata                      (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                             .writedata
		.onchip_memory2_0_s1_byteenable                     (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                             .byteenable
		.onchip_memory2_0_s1_chipselect                     (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                             .chipselect
		.onchip_memory2_0_s1_clken                          (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                             .clken
		.pll_lock_states_s1_address                         (mm_interconnect_0_pll_lock_states_s1_address),                //                           pll_lock_states_s1.address
		.pll_lock_states_s1_readdata                        (mm_interconnect_0_pll_lock_states_s1_readdata)                //                                             .readdata
	);

	c5g_housekeeping_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~rst_reset_n),                           // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~rst_reset_n),                       // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
