��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.yu�=�6`���؍�Â�"+�ˬ�`��`�Ev\�,�i~|~�����,k�A���;H�Ƴh��@�{9���k?�[{��<����?�FJ�Kb�o�J#��h��aR}֧0E�pP�'	J}�#Cܣ/�"�D���;b+���,)$����|�ű7�����Lu7o����JpYGǻsK��,��&�~�f����$Df�A��E�O29U�^�b��(m���8c��%g(M�|��_���E��F�㙅O�F8P#��
��s��Kə"���0`G"OZC�a-tA�' .�5������W|c=5�	;���-�>�*&�>��R�ru8���� �A����&��NWd��MQ��ZXm��e�T:ᤐ�'BUP�&L�y����)w��lÓ~s�l��ė�G՘�ЕQ{>I��X��/�[-�"5>B�j�駅϶���=U_a�R4Ǭ���+�z�%ʘ'�5�����O����,\����J�����~��>�5s��B��sp�,E�hӲAZ���s-o� ��A�&�H�u]N(������%��������[:�D�|�s�0��O�V�^�wkwA޹HN���Pe&&��&�?Qn";2��:
;ti�q�;��RB/%��KVT��gR.����F~9��XZNo��n���.}=��䌝 �0�K}O"����e6��g_��5i�۳=���CG��L��n����.M8Ix1�,��U�fPZq��e	�&v�;;E���6N�	���#bכ��Οh�!Jஶ?�Imq�q֢�Xik��o;j����g��D����x@��.�]IX	y3��X�3p6�?e��S��d�`V�H�%������Pd��r���޲�Q��D���&1���;��-�S��!�٧�A��8>z�^2�0�8��d�,�|FnZ�J���)���ߩs4�������[�F,�D�7!�@�R'��?G0IT��j>�楓�O�Ԫ�9�3��Lv������e���XE�py�	��WU/�n:l�V�"MXi�k2/<ơk$:T��G���������Ԓ�Oko'�ux������雰e�9P5�k��#�j��0}V�L�-�vp�T$�΢n_`S�hl�v��>�r&�;�2{Ƭ�r��hŤӟ���$*)���ȰЭ�V���-��;�<Q�Ha���[��3���;K��ܺ�-ZF��3e=��*o�OQ�	{Xn�4��R�s�({Ӥ���+�Gͽ ��ɪ�%�rcs����6U1����^�:�s�k"�`�R��M�j3삽^fp�!7α1�W��v�ҋ����g:��W�.����8��R����ı��nc��q���`w�b�%Խ6u,���tg�ڧT+CO�昊@�=Nk�v��֔�+�K�,N`J������A������ŪA��l��6��e�8&�]7���Ϟ�����7w=�[�co���t���Q]�P샬d�]�=�� ����R���'�0ǥg�E����w�+!��~X2�wz]]<�Z��jq@��=�h�(����-s�M�l򊰈��Ԙ���\	�S{��9��7���Cj	6�������߇�t����Et�j8,Da���L��ɺ��	z!h`����w�>j��m*V}"6�U�d��x�L�!��`���C1ZćJo�;�7�І;"�V�T�nI�K�@Ɉ]�ETj�N����۪G�� �x�饑�8�=����0��9
��Q���W��W[&?'�䅶�N��2��e���߫�ܟ��{���oL2��ǭ�ie�i�S�^��e1�R)�Jʨ)W�F+��~C1;�!�dDT�"��b3I��ۨ��7��
�Vu�;mC^�Օe�
�=����l	[O1�A��o����;�˥�{j�[B��|+T ;�@8\Ŭ�P��n�܆��@̇[@uux8X�Y).z���,�ڲ���C�c�n�mSz���)z�I �w�н��/��s���Ӫmpa������������߆hx �'�WR���>��Xd�5����|�VE�N�\'�X�� ���Rax.F۸a궤$��9^T��Z&f��Y��*x���?D�o`M�=�ܒ��KJd�y��y*(�����u��I�������o/���RTF:؆��z=OY�Y�gQ�j�95.���貮��R��*�>u%�gv��zo�b>7޵�
��c\XV/��� �4}���	�+�դS6*@Ώw�@?�̿%�љ�vـ��[|È�벋��m�+NN���6ɇ�yo
�b�Y��.�u{�.[E�nɏ��v�o�/_�Q�����*�ls핾{����|:r�ڵ�:�q�V����_���N���Oo�C��Fe�?���r%��L��U��K:_������d�U�о?�y���ٵ���zgF�(1�\��s'�S�ʖ�kF۾�'I:`�L�����1Pc��܁��z�@��׼�B�����.����i	.���Ӹ(�DT&�����R����ɟr�0BX��j���!~�*`�jG�|n����0�S����x�(��(س�]�j��V��H3h�N}]�$䁡	��4��������W/Ц�$�휨�2JC����XJ���-$�[i�(T5�ӕm|$.�q��km�K�t��0�%��UZ��0�����PIm��*�܋R��R�@�*��(eQZ��z,�4�����(6*'{����ߗ�wS��]�T:LgXNL=|7�6��k���!wNo	&� ��lkb���j۸Y� �bC-��a�2X-�ʞn>�a��"˻y��~�����i�u�j��Ĥ@�=<+:�d��'�1�g�e�!x.}��b[w��u��9��Q��Mz}2�X�Ìڟ� �Xyj��M��9үpEm�V	�vٌ��F��o��}Y�V>Gg�d)��r����iC��&�L�59�\˵���ۚ%_���4�s�0VF}�?����
D�m	� lC�X�S��� 
I��&0������-$�mU�*���E�öN��W�:��P��}�H&�HÖ��X9��mo���e�c��Z����r���}sظ�*��<���� fj�j!q�u\�P-i��V>:.`H��-�z�؏�y*s�ZX���#�,%d�h�UuB�Hj���2�z�������Y�tzIU� ;���U�f8F>9Owo�K}gXb1W�-��K����<_-T���d�L�KĄ����'�m�U�&�.��T��;E"����IU@ض��-�����u�}��:�{H�JH�fD&�w�,��������K#0��q�P�'K�h��3oP���H�;����i'^�G�\T"�Ω����F�R!b�;6�֑6�������~5���	:���|Z��\��ؿ���ڀ�]�_Jja���V@���l��ŘvF1�QjCqùv��xT�3��1P3}2:��q;HC���	α	��3�q�q�y%%�b���	���
�3C6�\�roV���`c�R�Q�sI,�ˣ�a�	"����b0"ްߩ���~���%�?qz�M��A	f�)\뽵#:����&i!|�� �߬�RzQ�m�k��D�R�<g�k��gu#�F��;�tzQq�!��Lr�J x�����?�]=>0��(��*�'��4US=�%W�Jxp����������'7K��O�q
�-̒��*��i����p���$���z�v�6À�N��p�Y�!��"�i��=T�P��O��b��a2�b��oJ��<'��Z�C�(���}�u�R�)-�e-(t��x�/��;D@vK:��=Ϝ�����6�!I�x����l�)SC�k5�<���x	��Y��!ቢ����g�	����u��k���i\�U{6yD�j�ݶ�ٷ6�5��ͨ}m�Y���R4�M~Ui��J>�ة�!�LT.�I��k$р �>���q��{ֈ�1�j��R��e:��k���P<�ʉ��d[:�h�J7���[��Ƨ�� �)�� �)���(����& `�F �������ualte��\b8d�n�9�i~1�@�i����nH/�e�0�8Ah��x�����F����V�7�w��(#WT����<���Q&f�+`�FGFø_,l3=�uj��k���iqF�ۻ�'�"���Da���Č>��ё��h5l����B{��r�Q;��+O���g��ԛ�kLC�7K��:�(��%����V*yM ��3<��:ns��	(Ki!�RpIZ}&�����0WČ&7�k:��I�]	���������
�c'�y!>/��Q_��I^�V��z�E5�<�j3��o��?���d��m�@�ҁ*��\�,@b|��:Ţv��`�ǁ�x�q^�zl?��K��'��nd�,�o��X�`����ڵ����ގ�wI�x�_�7���V��"���d�>>�!�Y, ������lv6*N�T\=��3þ������o'��N|3lQ
 v��A�*�W�O´$s�pRyr�v��S�.�`i/�j�i*>��aD ��tx�
�f
�?5�B�z^^�@`-�F�E3A��l���s�����1��W����B��<O��B���޴&L�@J�>7=��a&p0��/
(��Ǆ�%O.#xp؝.�MWq�蚠���U���K�F���T��@f��>����l+,f(c@���j>��쏒x���������pW������Ͷ����

���u���J�N��@�?;I��֩d%����̵�y�_�u���pB����H�9��Ð��&�艊B��y��5h_��}F��Sl�r�I'r�1ñ/����N3UP2PDϭ\U}����A�cyt�����8@����ruR���AxP0O������Βā��5�{1����rڣ�o)
�ޕ�����-�:P����
�'�V��<c��*�`��l��xC4��y��H�<�jN�V08�2 ����G��%i0Q�x,rWv������i���ҷ?S��l�h�A4$&�EqX�E��.'\4����Up=4�~�:N�#����.�
�����t�/o�6���]�[�T���H��qo>� 24������:e�,�1�E�뿱�)�".;@���n�������
���&F �7���������[ri�d��� �kCX_R���ˉv�4�}������yccsV֒t�0e�x��-�\�K'�zrۀאq������Ux�?�ZY�@��K�:WW#Y �o��3�c��RW?M6�8+���懸���I��ވ�����4�^|r��G����x gA&xI5�R�	��@����2,@������ΏD��o��{���`#�h K'q����(�ӓ�(�8 �ٻ5�v�x�8r���w�1��䔶g��.�W�������dv�q��Xg>y���T�v]C�����1�91Y���]�(ly���b�]����;���x6�#����.N�� 
�j��ʕA��16�O�ZaV������\g��ǹ�C�*tٻ۰x�)r�L$�_�1���B0�~��9W����&x�G�@��fZ��)��\�摊��(e�)1,@9�j�b���
kg2�+�3���e9_�..C!�K\��^���5��*=��R��c�t��"�^w�n�X�E�Tt#X̼2����D�+��H:�Y���|`�����ZQ$|^3�r�́sK[�I��[��5d��u-�R��u�@9v���=����r��~�\3b	��4AZ�V���&��V���*��#�u�[w�)�7��`��M��r�j@��ˣV���TK� �e���(��4i*�g��R�IHF�;U�~Z|��G093�a{it�;5��� ��~30\�qҢ�О
�!�>sS)�a�;�RMw6W���Nf�(K�٠�X��DGE��F �A[S�.��� 7��	������v�خ�Q�2�~�*�a�L)�X1�o���:L���J1�,.����	�5����������7W�_؈a�ĦE�j��e�5M=�G&wZ	�}mg�<��\�e!_�~녒��LpY�}_�����ƫ{��g�2���=�������-V$�V�����*�	�A��n�� ��r���]el�>?a�p��BpZ��&g!�Yѡ�èsF��)��zV
h[��
D�!s��Tf�(�6�%��#'z�A}�o������B&m��r(�Ii�A*m]32V�`~������ء�p��h��	�,SJQ��w@ ���1����&C~�lL=!l�[ߍ| M0d�+���~]z+1.�����9mGg�r�d��'[զ��Ӹqb2*�N��u����}Df��h5A�䌰���G��6���!�@�Z=pW 9�	߯\��� �ւ�G�i�9a���YO�����]1���䲕K�!\p\����t�����$bNM&�b�r����R�Hw~)�W�H��ؙ��� �Q�@��:��|�<���ܥ 4����i��7�;d�����b�v�]����aR$N���cY˘I)�K�pbc�[1�Ȧ���w�]]jni@ vŞtIMi�7��X4�?�X;�Пu��>S�D�r)�ˮ�X���[;4�<a������ ���������1��D����Z���<��-�o%y��f��~��򴹥ЃU�E��?��/=��B�?�[)~@�tUp�whL��;Ĳ�A#�(o�Ckv~~��w��m��/�-�����x�KȌQ>4��݂�O�Le������c�`�ŷv��b��K!	��c�t�C�[u�緑��z*ϝ�W�q�K��i�D�kѭr���8"��ɠ���Ꮸ`J�ʲf�o���j�u��!�N$rw����%�w�8�Z��������Q�:�-z%>���C?^(8��QK�H�{��\'wkz;�E�a*I��fJ�P��N:zF�L��z����5�Ch�u�й�^|.&�����_��]����2-���_0����� |8@n�X��=�����l ]'刡jUڻ�=�ԯG:8�ig���>��b�ˍ+M�oF�Nyx��l!'��BOS��L�*&p�p��Z�
�~�vEk���=_��嚍{�6����	g�� ¾�+W�
��D�����w���N�(�v_0G�Z"��σ�Q� ���6紤��%�C�LT�y:c鱄�x��	�Rß��LGf�1{J��e�)����%�8
-�����&��	%�4�Cm�ъ�Ӻ�����O���*��0�7�F�\~�Έ�M7E��.��mU|O�]߬Оu�[�P{n6,���K����p��hbPځGB�)�F�A%�4"h���>���-w�!y7��V�O�m |b�����!ApV��&3����N��i��Zӡ�No�8�]4�'��>5R/#&����f�:Y}������.�}~���h1/?fz�-�6)n@:ÂzbE��J�@����S�R�Pl��G�tvq%���󽏆S��F����늓M�70�s�ҳi&y7���)�a����@�_�0=e=4Kf�Y'�=q�ɜW��҆e�HC������ӡ�@��ɑxWzq��B4�ݖL�\Ö��+j����n[}F���(�X���X7�6��-vB��P��ٵk-E�2u��}�����=��!m�ȧ�F"|S��Ȫ��5n�!S���'M���l��ӺU�@wib���'Tt���g��a�|Ba[�o��W;|����Y*G�qЮ}��7>�Xˇ��b�K��j�I_tOt��{&��� +2wD^S(6b.�m���S�1o|��o���bܐv�p�.L��6벲 �Ib�T�Y]'�2�A���F�ߟ�~�t�.k��d��o��L�!�W�7�P��"S�v%�u��\<ݩ��	�d�V���O3IZ�ÖErw�*J з.l0/�Q�������b��y�?��4�+d5�!�V�F-OVA��f�E�LN�~���(��O��w�h ��.����`�^v�<�=�����{�@c��[���$����)�H��b��D��Pk����`��zإ���fu�ʷn��˙2�3#<u��.�� ���~��1<�{ @p���Cg(?��6�,����9���!Bh�}���
_�y�ؿ2h���uk��<h�^��B]��Q�++MoF��W�N�����0˹�G'�k!��O��������^ᴎ��+7j8�ƭ��7I%�����>ohr΅6tP�p�N���j:��m�{��N�۴t/��bx�r�)uH�g��;�}f�%�ߺ�(���f���'p�ko��v$J3-�f�~l�X�W:�֮��o�WR�V֞��
+d���a`�1�6"��&�t��]~<o�S�z d��מ��⦢jđڬ��>$�$��
������L}�ڹ-���Hn�B
��k�����|����b���O[<���3b��k��7�
��o-�~�ԅk�Cc�M �S�39�`���A��o�S_�ňU����"g\]���f���V��|#k���2k��F���R�7�Z����Y�����j�����(ŷ����#�����0��������}'~Hɥ�B\�un/��Up��Tw�Y.��*�{����(�kٖQ5���!cN����q".,;Y��-��Wq �������L[�,�@���	��Ls<����O{��`��C���� ���I�����L�U�c🀵���
��{�ГjR�j�$��TU}�afW�8�v�(�g8h�34���Vw�R\�L�� ��z
�d�
�o�edAC� S0/��<�T�Z��-%�i�Od��������:�bS��ʧ8��"g��ɻ�]j��Nw�h��?�] ��v�A����ߢp�f�?%�p~t믩���Uk�������y�{7���+�{y9sh���ʓ� �Kx]�Iſ��^�UN�b�� �y)<��r6���A��y�S&����u!��j���_Gx���86K�U(�����Dی�ё\���g���z�;�]��t��Z_�����I7ɔ��쨏������(fPY��)�:��)#:A�J+�Q�Vϊ6+����\W���G�z�ÄM(6����)�Ŭs̽K�Zʩ����8�xCb����{�-hU8���f���KSi.�������(��;I�nFn����!t�4�P�����ֺ�o)l�\��K�g��*�R�p�݈��p�'��Ւ�8�S��o���w�I������n���*�߀}VB�wz�@�O?
��&
̷����[}W��0���}�pz��4X<����-�u|PAv�<H)Lc��O�4��#J���Z��{�/5�d+�{<��[�}G-�m�1��$��n��
�dfx��dQB-~��~'I� ��W#Sć\z�g����p�s;�
��!.h6��!]�%4�(_w����<�N����ױ�-ߋ˳�f��|I�o,���I�-;��&J��4�jX]ð�0j]^�PDN�J8�����R��:�����.�R� 	���h�XM�N���{g���!����U�{���8/nMY�K �\6��D�"���5�YZ��L�����X3(��:�!Xo��[�u%9e��B�����M�{Y��G�͸X=��EP7YQ�XdXk�*�f|x#�������P$���7du�F�m��i��ރ��0�)���S�r��Z=�?=�I�l�C���#���̘<9 B;��`Y��C�b�6Th��L��E���_���h�����]y�T�����V���������_:��\�ͽ<!��u(:�y!h���Bǅ��IM&���*b������[����>���9��F��4���^|��"I=��,�Ы�e��P�c�����%����%�oh����c���q�����fe�-rQ�I��N�Țg"�n�9f�y-6����� XD��$�h�AA���*zR:���Ip�K9��S�IzI�ܻ�/�:�9�J۔'ѐ�߀���o�iT2�Ef�|�-ί5�t���|C�P~&*�|_~1�j(?t�0$0s�tI!���ns�B$a��*�}�g|΄������-���������/�>��?�r�C>7�j�DzQj8 �vy]���P)Os��"s�<*^��j�.(��Ӳq�#��{����󬍓���v��ThIH�&K���<c]G�0���
B5�«,tw��� $�N�Ǯ��C�g!E��d[�O4�r`���m�֫�^6j-��L<�3�s�
�pi)	���,�_.��9��F,�V;D	f�YX9�!�e�Cب�E����B��I'q��Q��T�
��py�c�9@+Ri���u��m�A���k�-��y�I�")P���Y )d��t[)�m`P�S������08/�s��g���.�=���خ�Н�,����B<��ъ2������y�K�����]�T� q��ޱ;��}u$���a��w�ЋI����*7���6�V�D7'D%{����s�8����-�����m69�y�9��糰���Y��¹y�!��/��������-���|$�<���V/�GmM��m�q{���]:�OVw�`OL� Ų��(-���C��NDEc���	�{��Ŭ�W�,��5rn�&����7��Ŕ�����̷�� IT��	%6�4:�V&�pSI�r���ۻA����JF�<�L�i�
$�"�W�/����%h/n"�/�Ƙ��X|tj��T݌�/�z�~@���Z)��TG�Hpr�1c���m[H�۠zXdҌ$�R�tR�@3"�A}���'�W�]�V�e>c��MC��\��9��W���an/��ݖt�Tee��IG�]N���g�jj/K���O��ݨ�<ĝ$�_�&����h��1GF�&����mtU��z�eE}�9x�����Z���5�D���+Q�
2W@ON�]����s����?�%���4��;�^Q�6�V^W�:��I�1��D�Yld�����/7'���x��O��aU2��	פ����4^��%���)��)�'�g�^���l�A$;녕���A����1�U��5I:���o僲�@N�+�5�ތ��Kv����fӳ��(6� �/W7��f�*��k?R��'\�\�A�c��^��]x��S�G��o�ׂ�d�DtH�3P��/�(&�cƹ�p���XH��N��.j�ޔb�*���h3	�
����0���i����ɷA��W��_&	�ϵn��О�K��
DU��e�q�Ɏ����j��E��Yy��H}�N�y�V�ί�a����(��Ob��Ato�B)��_�<�u�A����Ǧ�N�b^--�W��jD-=�Z�x�Z���[�|�C�ao�,����t�sF��`Z�jZ��H�S�O�L��"(Љ�kї�緲���@� �Ƿ�c0n�>�l8n0V3�Eظ�r/w�u���;8�T�P�"��C弻=����w�L�ذ��{�8�������1=�t�#i
 ��y�� �5;:@B��X$v����z��8�{м,�,��ړ��
�#���"!BO���mZ��DH�����Mڢ��S%w�PA���O��g��d�\w"��,N�h�jw�x����Ffˁ��+��ZS��D�����f�D#;^�����������:�d�#A/7�O	&@y=yd���v��N�sj���.�v�^��[�	����&7���;<�I g�E��ĪK8 �7�t/����F�*�?H�0M��.���_ַ�%�e>x���,ݲ�M5�ᯁU뒍ݺ��D��
Җ�q4��6K{�_e�m~�wBB��X��N��VECF�lr�ޭ�)�o�e�UH�)kL��xp�`�����Bmu����ˈp}qÝ�5V��������l�Ɖ�a��L�˟݂�
��*���2��奙笍�CVz�PE1QB��o�7@�"�/�7otB��;N`h~I��ai��g��tI�Z����r^.��!40������'6Pm�� �;`[�m�談'� 0�_=
�ʊi�d}�Nq25�F��[Fϋ�Cˠ|/�bq��&�cTc㆚-��l��%��3Oo6��Y���Ú<�Uq��%�>!�]�"p:v^�[m��3ts��4*X�,$gʱ��Y�o�W#1��3A��.SV�G �BNf.���]�>�,���=QL{�>i>Q1�鸢���j��Z&�U<R (:dE9""4yRGHƻ°I0�>����
��1������m��d�_Ǉ+4���o2�-�w��|�����@�q�J&�I��L���q$'�?S��GF������/�np 	� ������;���"���6x��am�h��z�k���].��������E��V�-�}w�����N29�K����^��+�C(A�[V���e������|�WD� �n��E;LȬ�!��Z�2���
��|�/Tو���e~'�!?������ֽ��hXɿ��N�!��yD�.�t$p�՟��4ĉ�����_5�
B=4 TZǌ7�k\zuA��z�lx�A�sݷ�����_k�G�{���z��>׀�Y�4z��_WLR���/����{�2Tɒ�٦j�u��y�ɒ��f{��"�y}+��n~�,�R��f��J3^�$�j#pN(rh|�(k�3�x��]�b�[��̟}��*=��(�y��1x�K6ё��p�U�|r謯�0Bh�[G��[�xC Q�~9�7��pX���^�Ky��*�Xv���f���7iK/S�id��r��#�i&>�m��j\o³���T�V�b��[-eӍ�4�nn</��/��h,�2��U��f����{ˉk'b��swg(g�V0�`�}��8�8\r�Q�E㼗(9������hd���.�_$>�d.���]G6��3{�S1�}�O ��,��͢�@���\�뾧��G(�I�d�H��� e�B9�Պ�ې����x�s��-��'`�{�{�:�џ�K�3��4��b�z��P�r�fQ�C�P�v�q�y^�W2>()W�F��w��翼�>kmQw.w���d�?���<	u{R��JYƐ��/@J�.�}�-�O��v~�0�H���9������p���u8�#�JS�����˼�ݥ�u�kV'�<Gް�����:~f�GzN�0�{A�b��AsX��xb>e-p�Y���1P�x�\�Y ɢ��r'���
	�g�>���T2��%I��<Z�߾~�O� ͊��p�ƻ?[��+�m;�rY�v�ĩ��7����+^��������3pi(%J�0?�z�����1������|/�Dr�J�fH���o�!q�Z��?���@wb��z��S�\	,F��rQ��!4	�Ƹ����E!��]�8�a�46�K3L�ljȠ����.C�	ƞ��T�[���Q;mF���}꘥`+))�J�Y:<!��pn�������� i�!��e*/�#�˺��l��!�I���J9U�%�HjB��#��p�fօT�������%�W��
�i�ߒ���(���X���~�G������F�]T�p��������9x_6}%��n=1���D��Q@]�<>C �oϲ6�QQ'V4�K�j�Y#D��̝^�^���7����+;��УC�w��:[5/��l����DW!��dL;Q���	�Bh�ɼ)����%��C%��P�̱2\1�ad-�C��~�Y>T\��wh��;/rE+�CgУ@��J��~R�DL��p��>N\�t���ي������w28=���I��;�"���u�G/7*O��;cLxd�����~ �g��C �	>j.�����1�>�T�-}�)<˞�;�s��b܀��mNw�cJ�/�x���ɱ�w��Z�����:ֿ����P�7���u�픩L�&H��q�Fr�!O�L�T��f�+ш��Uɨx�s)N%��Z%���/���
�:8+��	��Qa�� �-��:�b���;���[�o���Jf�t���7Ⱥp�S����XKZ\�`�ՠp��t���c�;�E�,f��[څ���ȉ9�l%2	�0�y�'�5��Q���
�_�X��
#����&F�I}�&ʉ���ojx�����L����O�Tړ�N;f���m	,�86�Xpg͢�7.�*ɫ�dOʽ�D���p��ߦ��ϘV�O=6�����	vU�p��o �	��dW��ǃ�Z��`S���=����w!G=��ּr2�:h�O�Om��-4����!۟��2��鵲�Sdߟ��*���\����]à���`�jx�6M��W�/�+�y@S:-�Z��Zat>�Zfx&?��C�#<kL�(�>�7�@Bz�������q`7�F�#�z������JSvs��e�S��&O''M�� e7���j�!��X;:G�ֽ=�/�}!m�bc	��L���x��W��/���ٗfI�akA�l�O��?^o y��)�UM�oN�/Z"���]���!�C���'?��1��䲙�qb��d���]�eGL�@B5SЍh!�D�o�#^B��\�內����Hw�4�}��/����8�]r8�w��o����m;G����QH��ʺ���X>fO�6r:��C&���i�0=�N/�,�@��ʮ��ec�4��� c��~��q����?!�5��]g	=�h4�fq#�mF�*�J�П��EzĮv-��T4�z�L¬>4�	7���V��\EE>I&��!U1Ij��L �(�R7{������z, ��`�"�)���2M�5
r07�RI2b����`���m%���ҶW� �0��sWJGԠG�\�b�	��퀽c0D�\<C��X.��iI~Tr~���	?\fkA���L��݄e��B�y�X��|T01Z�l��%��ww&q=U�4�ń1�m���F,��|8���:��]��b�KJ9��ъ�ܲ�k�0�g�v�T)wF��S�aV����fM����rwCD7]��˖�x30j�|��O1��d8?�};֭�n8;�]N�S䕻R�P�:Ȯ�X��?��J% f�c.�1MϞ4��-a��s֍��҅�_�d9�q�La��0�a+��d6���0�/����p�S��XOC�!��Ø\D��*�w_ܯ�̢�Z�����/S+h�+�0P.L��,Jy����Hsr�g��ĉ��F{��Ҡ=�p���K�o}�xNy�^���ɬ5�io�����h�'~JA��W�ۗgjY�o����W}��M&�w��GT�఼Ź:Y�����{�����x��lL�jB�b�^W�Sz�?�����w�us&Y��H���j�)������~�\�Ipw�IIO�̶�cDx���|֐)A#�b�S�I�b��ʫf�V'� �8IWq����9ڴ��aL�u3��X_A�tZ�/�C9����℘4=a��ߣ���]K	X � �˸� \U
%ds�#�S\�a���3�z�Q\�M�T��p�I������\�;Q�y E�p��D�FI�䛯��pʶ�q~��]|�V��)�i�I��x�>�~r�2��G$㼼a�5��q���C�jrFR��ۯߑ�GJC��MHQ��g�,D�Hww[���B��Ӓ_�C~	��ĵ$�j$ke�!G��T8tD�٘���.���#Y9�$�¼�V?�G6�7ȶ������K�[�ɠ��v����=#�_m6��C֕�pɠ������T𪅯����"��q2� L�A���%���bÎP����fG�����)dl=�+�JO0M-�rZc�>�]S�N�ߗ?Y�����Z����b����_m���ݗ;HX_./Q��X���V�����a��k�)7��X�0P]��5h��lP�G-�uW�?��A�fk�d9dU�X	�Z ,L5)j]���a.���IA�K�릧���Q�Y	Bf����J���`���7�4a�;}���O��آ�곋QR�� 	;�vp���@_/�Z[NʱceF�3�HdI����ku�A,���[��nz�������~���/u�f�M�41�t����������&C�m&���e�2*�7�r�3D'��%�-f��P�4?	�,�]�����@�$�v�!�d�F)t��ĸk�J��ގM�!Q�?z�*�!i�V����!u�AK��P ����]!})��!@.8C��{�Ϧr�A�z��kz��:}�K��ča�h��	.��-��q�V9� *���0�T7Հ�vF������ ̟@"3�v�!t��1���o�p�V�[ߘ9$ۘ���V:��U9%�0Q��&��"�g�Fh�{�WU��3�`��-�}��Z��1�#�Q���PB�f�BkB#��
O���o&4�֜�ݞ���|).�7��X�:�ٚ8�gY`�2��զ�ER�l�HM�Q��=�:vApag@{Ô.)㉆�Q.p�"�r��[9�o&��¥A���zJ�7ujT�HB�s�cE���)'{���p��&Z�B9�o�=�| �LN�!D�Z3�;H+n`�+�:<1쏥;�;����:�LZ�w(TAq2��ũ�\r��W�W�rSq���o�*q�	�-ƹ%BM�d5����~ft}�-9*�`Wƣ/�G0x�C�0�Uk׳� ��j�2R�0�u�o�����D�|'+v����;��I�"	Y���jωQ��Fliy�\���s8Yd�S���*I�hŤ�$׵N֦�yF�2��Y�W��e��p|�91���r����P58u�߮Ά"�>��uwq�h�<�Wg��>��4��s]:;f��NhU���/�9�Vܻ���*2�!\�I/*� �������
$�)�:+x'��eP%R��ת$�D_	m=Y�J������f~��U4
K<+}��Or=��c��3����x��8��<����w���@�Yt��@m@�cfR#���Ш�T[r~�dʂ�{-tڇO�u�Cq�C�O̐�l��/^��WfYG��g��e��R׃R`�����?�3�&�u�ڦ�0^�Ѵh -J�r��������.pÅφ�V��7�B�~������"�zx����|������w���N�ݮ]&5ݩH�i1��Y��5�{M̽����b�ʵ���>?&x��1 ��wp��x��G�_cz���@r�������|�0��?P�����?��
��xZ
�}M�+�_��^��|\�������eϣoTm�*Z9��p��	-[_E�2���i�X�-��KW�U�Ak-�%ͺ}q������~2�Nq�
�7�̠�r��q6bk
�~4^��`�+����ߔݵ��/�,��iqH*�;� [E�&��"ޑad�a�i�
f�B^�xn:�E˵
�32t��qx�
��ЍF�O�h�~^I�Q�e�P3���4�Ϩ,H���C��Ӡ��D���9CěO�-<$�e<{R�����F��%E;j���2SI�����0n(f�k�C�+�=#+�[~����P_����,g�X������ё���LE��k�U�����C�7�*]�Cx�l7���[�Z4���W|.�������.�J����%8��0c��Ω��!6������7F�jnx=�_%t�x��������qrd'\���x��QX5��]�y��]���$����{� ?O���}V�����Z:٤a=��6L��+���O�S"�� q���h�	���i�<RLe�D#96lE#���vy��R���"J��_�ڽ���^�t�˩�j�.a�H���B��N��P���-u�G��|e�GW�&[��8�/y�?+y�6�$R�!V�4A�'ibHm����颫�{�!<�w�@�_��w��,Tj~x|�������ֲ^�}�\x��Қ��7
��l45 i����0kO�zw�� �Xs[�Qd�u��6���Kƪ7j�}R>a��-,i��]�L��R�����K�K7L��O�`�`gQC���Qo�����O�QD�HKPC����5UuD�@۴�q٦�����ǾĀ�S���L��/�*�8��w"�02�@pH���CY�u*�&�k����3@ �<[M���&���\��RtR���D�p�)%�2toَ��^�Yd8����m�X���n������OE!�W�fD%;��mP�;o���p0�6b��_�a�i��hۆ;f_B�;�H$��P��V"Eqէu�bOVD�頻�RW25b��:9Z����,\:wё{���è�a2��3(�ca�J����&Y�V���'M9zg���ǵ�c[�m�K��2�"k`� Z$�{�鳱�ތo$O<X<�f=��������2r����u=�w�d(�}u�WMj��P��魠ј�I��o�{'��p��c�0�����'�$ݍ�C�r�}� 7���C�{{,w{J/�*d��f������3$9H�Y���$�^��c�I�q�X�ҡ�I�I�K�.�=�����jch-�)P���N��0��W��|�yJ���<Q��⣟n�K8/�(�5��HS���hmk
�ؾ�5_CZe�?Ⱥ׃��G���<�p�C��k�v'O�����Rۂ�5U�יE�/�	��1OZr�2���՜,�ە���t�MmI�8tmg�2���=VD�L;�I�S��9^���%Uҽ#�*<w3l�BW��R n�`V� �&@�>`@2� L�">��~1��,f�4��!x�ֳ��<jH00�- f]�L��T�����`uA��5���$�*ŉKߡ��Vf8A���j�Q��7;����D�S�D�7=ܣУ���D, �m�+�u5gz-cbG��ps���s:Q�5����Bi�]fAH�� |>O~�#�Ő@1��iX'cZ�!ح�ۊ"�9�H�<��o�[ >gg�G�z����W@?�H���	��yJ�W&med[WE4smw�x��pyAA��dS����z�8cT����?��1 ����[`�N���^�n7Q=�D�9sS0:8L5��C�tg��ο�X;/�i�!�5���(V��g-�C'���x'��k2�V���n�eunͣC�L�EZI��^�$o%����
�;�nAR5���ˁ� ��+F`��(����2ࢾ�a�,K���q�3���}>ǰ5��ą�c����I�y�lS~Ǜ;����Z�п|��y]�V��b�B�۠�Þ��2�Z�H^�1����k�r�T��v��1r����O���JW�'����b+�j���}~�����u)I��
�	y��=?o[�ʹ���"��~�?�j0��?"�������[��B��K��E��,���ZB�DL�H��a^��T�
�m
�k�p�������f?�e�1�ZY�yΐ��K���T�_d�U�B����7j��D*�C)Q���
�	�9����;tƱ��N�3�Gӵ�~�����EX��Zωu��~4���J�!m���iD(ߟ�a��S&˂��F���{��q\T\��f��G���)$Ȟ�?�S���Q�E��|������uئ��n�	�m��<�#�6,�*��?�|�%�������)��1����4Ѝ%B��+8	k�i�<��ݖ���<�۵�9�De/���H��P��*:�%O�g9�/q���^Z��Aj��1�1+½�������޳u�֍[����8}��e�*���� �1��TmC�U�n�QڀBP����}�qc=���鋺��.@������ax��Мa�.��i#�ȳ�C_�a{�ãH��[Eڬ;������6�2{��9�Ҋ�omՅ@D��d�z>�SZ5�и��XX`#4l9��GN]���h��L��Y#�l�K�t�N�<�?77�	6BAO��K��X
�ӭ�s�����H�/��,�Xb�d��q����9� 0�bvCu/M�֨��Q�!;.��C)S�$� �x����2�[�n瞂�S7��_x��9ض??
�ylw5��\��А�)j��4��==D�=�%��oଌ�`�*�r�&(���c8?z�à[���R���?�I�����щ���0��&�B>�Ȝu�%#}Dϓ������k�>1>�A�� <	�1~d����o�m�A��L�o,�H�*�b�4Z�qV�Ђn+��	��f,���Ĥ�}�S��\<6�߂��6r�F�ܾ���}���C?A�'�閦tA�L�m���bc���BI��ķ��1�����oX�#+?�,&�!�o|�uPL�oA)��18���7�!�I�9�UM��.�}�|�FƂSͦ�v@�����:B~�)�����I�ե�5+C�g�l<���kgp���v�ۓ_�(+�R���N��'�$V��a�~/�h�0Wn�J������~��60�Sp?39�(��haUn��*�T�-��w͊�|(T�9a�kܫ���[M�|��q8���q�I��h���;���W�
s:˄	�]Ċ)E�9B2�vt��Nɼ��?��ƹC����תR4M��pFhD5߇ѓHq�'��LJj���	zSɌ������DĉF$և��k���C.�.Q�Բ��|U�%<�@K�[�23I>v���V=-��:oS�Ԋ<*)^ҙ1UD�&����׮Ƙ�r^tGCeӥ"+U���1�Xʂ�Is�����qv.b0��d4���7&gh�-���x���gȁ'�*N�"Ĥ5����P����:���;����`%��s���O����'g�g�����T:�"I��3�H�"WR��i=�1�*6J�W�J>�q�!�ϗ����4Ҩ��T�M��B�z"� x��Z����%,QDmv�b���
�9+;�.%s��*�9�:i���&�
J�|ڭ�wD�k$	�;6�*Z��s,���	�rh3��8��c�q�,p#��Ζk�4��$?6:΀��G8��-M���.�)�p��}lp�@�6[��ܝ�5o� .����a�[���Iglh� ���GPϏ<�;J�
�^�u75�����l]]���쥀T2�K�����s��E�ж	�u@9EhEᫎ<�F<���LB߱D*Dz�	v;�,��0���嗛G�(��䶤��r�2:|vb>|H�C�Jq����߷�C7l�u�΢"@s���Jv�ҟce���E�t��~�,�Lƕ�����"GcC"�~�?�ȍ��g����s_������hW��Ꟶ��`T|R�!9
�an���!�.���(�9is6Kl��)��U$�����.*��Ge��vF�T�*i�?]�cڀ�|��¹�$U.r;.�ŠiN�*�����u��r���X5�����jEcSH�+z�ڱ
��w���{��h�K�K���e�	��yE�K��+�rŞB�@A
���2�}�0o$����x.���+MA"�,I��i[�l�q07S%R<����(I4I0 g�۟�a3�s)���u%I�ޝ��(����ל���2a���L�-�&�}�|܁'~|k�H�}��Z�F�\��D}# q�"�p�s�{�$�2<OR)�.4�x�q�jxs�ф���
�v�*sEu�-T�!D�Ԣ�D"�P_���ϵ� �h�ͽؗ��n�	��#)�2L��G��|���>�dm J�G�l���l[	P��$Ei5��ݫ�A�j�?]�bx��([.���V]���^�fn�A�,��� �S�Q�5��-nD��T8�d�T��:Z�hf5����&�ǔ�|��;��`hc�`�j��ź�s(��p���L���ې_ǰ�� t���k�ܟ�~D|2��[M�hx⪢��H�r��E�◧, �?�3�?;���5�p6�#L�g<���v��:�Wɓ�Y����P�w�`�g��;3��!�ԮS��{`�l{���Z��&gH��eǞ��_��kw��)�q���N<l�������c߭м�pͫǔ�
[��iDy�p�e 8~ʩ������i!���8�#%yn毢��Oo�Z��e�ܲ��ʤ��O���/�|�~pm�.�)�6gNZ�T쪹��n`�y8kQx5�l6r`-h�94�{��
�vI5fR�-,�`�B���R�f3tNU�nZ���Ձ��~5���!��;ヰq^[�BvTz�_�a��l�^�&܁������7�i���z��p/�ߨ�9l���J��WX�(��&�E�9�7������o����,�([s�T��m��Q�/�E^\�EH\���:�<f��N��P���t�h��ȁr�k�Q�N�V�mnR����h:���͡�:W��aě�{�wv���oc�V�?�/�� 1�s�P���Hʨ+�PlXEi?n� ���]..�ʅ��?+�8��!m.��`��I}m$D':y�(�oA��1_��&�1��aڄn�����r#�b�:��ZU�z^Ӝ�ϗ�%o8%�+:�Q���?W�2\�|�K/�Y��b��kăi:ua���F �z]�g���`;��p��)K�9�*��Id��5s����|"T�yM5+˛g�
�}g�����,��D
5./���Ѡ0�b7:]+\.�
����
;��`$&�_G�#>�j�k�&{�9��TZdǶ8qG�T8@�^զ�ٟn�p�.�yG-C�� ?���d��N�(��H-����[���k��og@;��D&9a�%�wH�~�)F�o������Y,�=f�CCV
WF�����������XG�oV ]�~?�m��f���M���8]bm�5�Y���$�;{����MpIݧ��c�{�J/�Aվn�w���s�hK2���ӫ�H��hrFwZ�6��Ċ�UL��O&ЅX�& q$��A�����+�����; ���{��5�NT�����m���}���c!�X��L%��.4+��ƕyr0�g���3����0��0�[����K���iڂ&�7[��Vp�;.�w�o+E�O�t�U*��N=��J�����E ��X�(IJ��	�87����J tJ`�0�D�Y�S/�^�"5,.0����V�tc��T������&e�c�渌�7M���a���
��ۯf%���q��"�H;���YU(V���p���r�~
���)���}�L�77�<o��с��M2��8jyH�y�Ǆs��J�Gg�Q��;�������� u��a_��[��)��Y���?2@ Ϙ��+[%��7ɷ}�cC��9�M�{��V�y?DfY�~S�f�ǭ�+��'~K@�\���u(��G���=$U��^`�:9�ίS��:8�g#RB㼏�=\�N��h���bU��U6nn:�����uK�^��q����|R��v�)���Up��{l#/(��`g�kz����A�`j ٺ���Pڇ�V��un2�9g��x+`��5h �
-+����|Sk�G�.9v�n>Փӑ\7`πn�Z_ֆ�9�Y#&͒V$�' Så�A�7���^N��=,DnFB�73z�np�c�.*�������u��s�E������KIA'�1t��M��t��`z�OG�"왿�*��,���\/��U�C�Z���^�����o�8�zm���b~&]��=9�@���)6��"����9Ւ�'���u��X�~>�+�w,d߯���mVb���T����ФG�eT�-��<�����>l�g�e������T��h�g���m��i�{�ߍ9��b��ff����&�".���v~2�����Q4,N}�)O���{��I7���1��ؒC!v�pr�5Mfx_�>�F-�
4Ի����� n�$���>Tޑ�������*i;_���
�P����m��T?�{uMGF�q�r�Z�V����k<e�e���H�s�@;�܄��?�e�K��g�:�.���,��̃�,�
�A;�9`gh����Vߊ�%� ���I����",]!n2�Z�`�9mΎ7P;�F�����5v��w��p!�(`�� ]���'Z+�S�ٗ���\)r�$�(����
�#����W3?_7FNE���⑈;jN�4��YT����k����T|c�$����qmAs��i�����~?�fbq�Nh3#�Ba4x���a�u՞�|��6�d�_���R�'�?��dC,N�y��o��v�ܤg����^��*W� 	�Pa��\�_�No�;��(�3QU;�J�"[��#8JВW��&CH;]2��k�T<�V��2˧p�*�*������\�R��9�7󊉘s�g%w�D�C��S�N�◒װ鯴ZWcf�g�q���x~�=^����7E0�۠����چɻ�����@�]S��t&����C�/��p~��OQ���[ ����<N�kSPFX]8�I"�>1��`K�c�&P�*���mÑ6#�6���Pi�q���{��#KQM[�a�쭆Z�+��V�I9N"��Ģ�	8;]�!�/B����./b��$�R����Mv�m���>�#��D\�t]��,��tZ�M�,7_j�F-�^B1�SG}W���{V=5өIpTI��K�w��΃�`�?���Q x���<����Pl\q�|�Q��6\T�-#!�թo8,�x_Og���#\%'�@n�8��6\�:��œ���-��A"��Š�vɀ0�r������W��Tw�4�IRm�b�@.���;�o�R �뱫�$����KV���mS����7�P�ڄ��ű^�n'���d�ΰKW{ğ�C
ѿ�3r���aX!�z�<u~)�]���)
u�ĥ����~�S׽o����坿 �v|z�s��?x���s룫��g(u�I2 -%<�r�� pf~L �o7{kJ�d�[�6���(����u�h��Skm\B��v� *Y,��LZ���<^�(�3(|y�"{��bF9�)n����#�H~�۵ha@����U���'(�.u�&�,��N_c��'v�R��-�E�uk'b���w��U��)��$߄e�(����U���2��~���Hs����s?�6��_�`�\/r�|�P�'����*�=?_�t4O���3���ġ�332��^��}�,4��q����s��q,67���m��Mp��;�����4-�f�����,U2����1z�� �e8Gv���tSڑ`gJSi���Cd��.��(ZPX�(W|Hz8w��?`��ǚ�y[�ɡ(N��O@}��W��K�!���B:�t�f霽����*&��>p����^��N��̀&�b	�/|��B��m����5������{��y�IA�>�h�VK�T�����y�z���:2�j�i��٫�D0��Q*̭C��\�}�|��%V��� '�y'1��9�u>�x�����}ڏ��.ԋ���B\��'�9���ߦ����vE�B�)��OW˯S7�!a�.�a�?Y�C-�Pܓ�O���Q��)Wb<cb�]$Uj������#gYJzƽ� xѮ�		�R�/ y3SP��1�o�t�#R#h�P�� 8��H�S!ң���`J�.�C��D8~���n㰰�Rv�YZ���fݧj����3��M��Ңy�ĦK'�U��}�1��N4���Uk�C��
%���OQ��et�ӹl�LE�V�/�XbO����9�'B�v�e��~�sq0���
��p��d㍅&2E�GpV�	��V�I��mS��t����*=ZDKR�u).�0rwDm�Ф��(�,g��5� Aq��]�Q)K�B��G����-tW���1�����Q�7�U<��i��
�M��O�{��셬�����Í�!7ژ�m�J�w�;�U̺Kw��.��l���x��x�؏=�+�5���?t#�IZHH�󞸎����?p�m�Uf�̍b�퉂���1R�Ҝ��=�
q��ȹ�N�����^�_#���ki9f.��.�����|<�sZx�u�y0;:ޓKK�����&��f,�:I�⭍��Y�02´�I�
��'���»�C18��\�!i���0��s�� S���r��k�*0DN�'�.��h�VI�pS=h�eM�"b�I�Mse�YO^�g�F�Xz��=�ý������!W�"8�ڽ����Ee;zGY�������D�?:�����j,d�	���>�>o��f(�"���D��+=�h���U�ԙÞ]��1�+�Ϙ5F���L�<�$,��o~4`8�W0�bۻ���\<m�kN��D��J���f���IB��K���IZ

i{%������NXg����tN���(k5���,�6薔H�HP�w[߽4���^����� _�V���u�T8�v5a;u���v^��p�p*x��`e�2ߢԤ�����>f����F� ��Ld�!�,]_`o��j(��[A�|.��HM3�K�ξ�޼=e�ڊ�!'�,�X�x�sʽ�X�rSb�����Qj�g�	$f�lE���_�l?�h��,^��iwH�)g3}`q;�y/��J�L4�$�`�S�F,\���s�
`�H�k(����8��Y�֬�m�ƣ��HO�rrߙ�Rq
}EN��M`gq��Ĭ��[}
�>����C�x�?`��a�c���Rs!�8�L?K��V6�3x�R&\<��K��<����%R�N��Pcl4d#M������͋�s�U%���Is^x}���S�l��ҵ�9Ϣ�o�D���W���2br��{2�q��ů���u_8d]�©�%���U�Yw��uȩ��y�+1��QKre2T�~w�:��@��J�PU!��<��s"W`o.�Ƨ�R�W�n�6���� =.�v<�	ky�NUB�PB8�!o�ʕ�[=E�'�X�δ&Q�xD�@�Ub[��U�s>L6��t��l.	2� у�\+ڡ��fY�賗��n8g��M5"�Rۋ����J�Jy:�vw����S���V\-�RZ����� �v�&LTj�I�i)x�Qv�q���r�,<�:���B��L=������>���>p����Ԗ8$7ZDI.N���*����Љ�̳~��o�N|�-��p]�|�5���l���j��H9s� ����V�١���les?m�
P����ٷ�UܬN�D�����-�-�ˑF)@y���|S�ށ��*�=ߡd�8A�uS9��W��J�^PP��wv{X�ׇ �/rR�ZP� v��_�x�@S?#��1]A�3�ٍ��A�vju����dT'i#������g���{��t���\W��ɪ�V>xF�+(8�� ��g �xQ$0"��@.��<��AJR�띥��P_����cs�����7/�1����X3R!����QDSEZs*#	�	Ta�r0�/�W��b"�Z�O�g5ڦMk����ҞN����i��j�;���h�}���k���ܸ�<z~.u<B�6F�A�5eI��c�Ż]w�8��l�uw�d�4���mC|Rr���(׃��~�D^�8����Zw��߇y)/,��*&G�u����+8; �{�J�Q`9��5C�4���$-�6,�ل�=�Ƿ>Aa
AKt�<ŉ5[(N��'�O�j�*j9�|�fˣ gbb�zB����R�-D�Ȁ�ik��w!x�2Ţ��X2��Yo?3�X�����������uޛ�8������?p�&����(��s89�T�w%�f��L�feH�t��˙}����3}��vRP6Ɓ��.����S��\awm9#Ҙ�������~�;̄4�&j"����>�7<��Wq�����q{�"�	�v�49����P���^�P�*�@�k��Tp�@���F�Q$��xBj�QXk���N�H~������-�2�.�U5˧8�<�ͮfC1�ca��-8i���͸,��:�y�,��Hd��۹�gD�;(��:�ԈD�ds�G�M�F)J{\8�r��dT�=,&uN��z�y3u���J9��ӊL,��Pݛ�Y1�tC���	ӒU�����R�,g��:�D��-G$���*Qe�5u�,;��el�2ݡ�aL�В,"���>�Z��y'�o0�X�X�l�q��p\?U���LϹ�����R���B���W���5��7S���'�����F�� D9F?Ƌ4}�[�,�p��ߛ:�k.3饺��O�����l�.�'�-D�1���0Py��@{+lZ?EC�Wdd���� �����e�9��^D�ԭ�Ss�y�}L#�'DK���iJ��u<�TY}�����[����/��w�茒8_�Ȕ�P��Yaq@G��8���«�a藷�o��w�t�Cf�]:R�6��w�#�v%��1Շ���$��]��N�>���Mr�Ҙ&��\d
g}"# �a��� ȴf���4P��o����mN���ُ��A�٩q,!�&v��=߳}�j�¦�CB���Wrc]����Q]���~͓��Of��a�\��3��\��=¶8S�PL��c�ą��L��q��>=Ǣ�'�*��8�U�
)Rq\o�1��� .D�t�JQ����V�eg����Vy&��x?��%l+�����d�i�C�X#{ǒ��\J�T7��;��"��T�p�����SB�K���`�[�=O��z��C�2�[,᰼�N��"b3�#�$�0ǩ���T��J�ϕ`p��E���!R�^���
��6Y[gB�P4� �`�����6}#��D+�u��yOcH=�g	��t+��dr��6t]!s��Q�w��Y�ų�VZ�\O,���܄Q�:�"@��i�����#���<9�c����L��q�MA�^����OZ"C���Z{�׎��B��N�i�<&�ZQ���L5-��D8���j�>��R� z�0悞7���`[�{�G��&,a���0�"ɫŬ&^�}������RV ��D�5<�_癭�������"�k��`%oŏ��ym+���|Q���%�.=V~� S�ڕޛU�0��MHlp+ � m3.o��k{�#�f����B�������1	���3쫎t�%�?Z)�v�hid;Ж*��"!�X���F�ͺ���U����׳j���-_=���`������Y��n��&����W4���H/Y���f�^K�	�Y�.׊�ҁ}��q� ��_�s��*ӽ�ą�Ay���F#�֢Ŏ�;ṫ��k�{$����=���{���,��HI?LJ�2�VT?��E�/o��, �]([�ȺH��|t :�Ⲉ��6a���d��MYw�1^B��>������Z�ʪ��v�@ե�%���W��6�R��$!2͢H�͛����\����B�X�m"�#e5�j�3��#L�N��[�>`�4-`
�Vęڌ�	$�C(���8��Up��r����e5�>e�,T���g�)zi|�T帻fߣ�o����\�JSg��Ɵ�_��R�����k��Uh���'�`���\Z�V��I�eVB8�.O��n��y����l����^��W���	�?���0�]�e�];du}sZ