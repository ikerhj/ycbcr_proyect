��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.8�Koꃦhpu�Ű��"q2Ip���$�f���d:%,������yxc�9��a�_aC��k����'����0x���aIP�C"�Q/$_��-��ON����Y}�g��b�%���7��IsI�y�G�7�'2��h�	��sM��Wńx��n��Ög���	kK5Lt���j6m\�8�A^T��*��&�^��ݟ���_8��"���bq#���@��������x����L�jJ�%��ݼ�N7и�X���c8��e�ڱ�W?��	���V5D~�� N,�@�!�I��U$CQ��e����8��q�u���t/�>`r�0���O�hs3��۴�_l�8?����Y��F���u6k@D\d�Y�$|�#̦�g��&̤sWDm#J{��k/�ʛ�=���/R�i�Ǟ-�2��x�|����[3��P��R�K���d�����F t��N,*�ג��k:3g��[�w�dy6oc�
�y��0mȠ�O��cO�`.�e^_{�!Rb�r�t5����fE$1U������2�k�޽�$[(���FB�<ݫ��d�}.L�u��Ƿ���]f����	K,��`���J�j�^/r�|zC���#�W�;��|[�z�S�E"?w�����#w�1��M�bV)�rTw��#�Q�s�Luy��M�7�j�Q?"��@�A�~V�VL���uvF�UP�¾��ឍ�2 ձˤ^RhՂ�vP�}U@����0�:�c|.Ϛ�_�����\j�(1%��L_��4�e/�PN�#,����5�M�y�d!���!����i8���JނL�1�4\��/�M$(�
���s)������뙄e)'%�7���P�)<#��y� Hj�sK8��1�e1��"�!��Ja<=B\�����1�v�ͭ:�����we����7�ҧ[�j�L���+i�SDo�v�z��C����Hc���p�d�ָ��Jh�X7�.���3K�9�8��nQ���Q�dpU�k�l�!m��Q ?�̀��Up�C�^>�51�{����;\�"���W✍��kq����^�YGnOذ�}N����l<���[�u�R�'�(�LY#�¸�t_xz3<KUgt���0��={U}G�Nv�?�3t��e�/�v��j�+O3}��k"n�y����X!�?����ђ��s�?�8jOՀ="IP�e_ f�Lݘ�w(��@R�#�)�)"�,_8���Ք��T����/��s
�;��2~`"/?�y���ܻZ�}�<P��%���_�9&�>	����AA��bQj���\<p�Z�������I?e&��z�����8KՁ�^XK���'�'�s��#�[�N2&+i�T�'��2�ގN�R��#<9��GZ�����o����*�p%<	$�6�?v��4��C+pRjv�g����tQ���)_c�Ӓ�%�_j��k05�V��5ڧ��4�2��ߜ��E9�=��P�q�w����s�{�g�~�H> X�;�J ~΀�Y���p��P�+EO�8��5�|D� bAI�2�)H^,{ �O��V������$��R��z�cG@'�}18L����nqu���|tb#c �L���h�N6�ú���%��')��{�����p��U-��X���}W�I�\��40 ��K��;��������l�B�(��1F�t�͛zGS���K����xl�hz!��xL<q]�\+�AH��D �6��t?OD�!��Fz�.� y.L� �U(�X�C�]
���p_���n��Ղ)+c�z?�e����* ��|�ҁ���V��B�H�M��t=�ko���Ӛz����b���c���\T�SU7].�t=�8���b��@霳䐱tl�A_�)��dm�������|Q�I��e%4va5`��.�Rsn��w�C~�ް��<bi�5��c�G�Muw8�YW!����9��0*����CjX��-@��� �7��`�p��]�P������գ��\n�����;��i%�ӽ�X�^K��F�U�e@�]�������Ef4X�)cbbaG~���P�"#�X���$��e�i�Wn�^T#61�>���q!��i#��8ۿA��VC�^ӪVN붃����jg�3UcA�?��S��1�󷸨p�?��a�t*��!5c/r�*�g�=m��K�H�n�͗7q.�\V���`#��)`b�2Jj_����L��Յ��MZ()��(V�]^*s�eL�t^W/V5)�K幨��EK�9}z�9ۍ����=L���-�w^RHqJ��`�)�-^
W��� ���q=��I��%����I'�����U��P�`�9��U�)���m.iy�����0O�8%ŲQ�L�~r��W+�r��K�bl�)1�_���"��a����"�F�c�L=��l͉���)�x���{��$�����6ʑ|!� �ڛjJ�6���ATUE�.�J�+z��#/�5��z�}�0�q���:�4�F�"6~�b;R�ReF��<���x���M�"e&A��.��;Q�^��2x�^�Y~�fV��Y����tF��k�O_�L��5[l�c~M��% ����Qm�}���.���1�1@\�� p�7$�\�[�-خ�+fﴢ����[��9z��<��R�"(+�!�?	|[ �ֵ�B��`��^��k��\$�1��� ��p������$ ��w=�#a~�v�P�d63+���s�:�5��q�b���O&y���fΜ��D��Q�3c�~\�9e
Ђ�J፧����otϮeAM6�E:���f�5('��M��R>����>\n���������#\Q��K=���:x���²n�*�t��o}	��1�^^�g&�h��A]�v�Ek~] x�s�� ,��,@�-����.�&i�b� 4�b&BG75aI`���Σ���A�X.���dF=��3FC6#y
�r}RlS�>(�x'NQ�F��d�)ȼ�"�̋���Y�eB0>96�R�N��r5�ʟ.ۖK9"	�l��Ri���NN�+�/�j���� m����/��w��!�q|A!��lR�g"?�8���f�`yw���k�N~�kC5O�Е&=��j~$ a`E�H�V���缘��gz>'ک�~U�	"j۔�/$�.���H7� �\ȥ����wv��g�n��WX'�J�GC��x8'Q@�l�4,�P��%���}���q5#7I(�4�$�W�Ԩ��d�yB����.)���W��Yv��JJ,Ez�#cƀ7+D��S<i�S�D��Z�,�=����Oxܤ)��L���fa�&y�k3�^է֚F)S�y���ηȒ�^�'��r*���fA ��ذp~oy��R\R^���Y�#3ox�܍nȊ��/����")�eeF�W�H&qf#yrY�[rS�.����%fc)'l����1B����� �o��![A0��5w%u�k�*&	�ʟ@"���KPV�y��g�C�ak���Ԃ�����h6b�[pS���� j�����?yKSz6&��Mq%!|r�d������5 �BoY�*��H���'�2Rԣ0mx=!U���8�w��^u��P�I2H�s�BiE`�T��7��S�reE �-�j��L�PX��Ʈ��~>B6��!�����:8;?F�3�#� 3�O�؏�-4V�)�,_�b.�J�hNU\[Z'���B�~RF�9����Q������C�&�܇v��R{��r�K�6���-�ק}�%W˷)Ɓ�e��J���y�)�)j�1�i�_x�쵕ث�:���+Y:��.+`>��6��`����� Y��V�A�Z��1s�tOL{��R�~l�n�6���c�����I��0n&R���%"��ZЁ���g
��|*�{����Wi��Ao,�s��NWWR�-�l�=M� 6�q������Ӹ���S�&gm)�O[{�~�q��|@�41~{�t�H��G��b��V
/�n�D�p��'6=�v,��:;?Qev�Z$��b��]�l�=e8��I�L�q�9���2
/ V�WVp
��s���yŠ�V軃ߤ�Q�F �{S���@s �Ҵrng{���~�7|�fz�Zݩ֌���'�)���i�#��J�Nϐ̓PhΨ<���:���r� ��=�?��m�S��i�T�J�0�EF?3�@� ���Mt��w�����J��Y<�e��C��ir/�� ]A�Ӈ�	ȅ1�������H�m�~�� ����>�#-��M�Lui�j�1��+�ׄ�:Xw�D�϶"��R�ȩ���ã������"9%��5.yE��t��w?������=�:6�Kt�_�����TE�~1e)�?i�%���X4
L�]�u2 ���`	X�]:G{)����?s3k��Ua�I�dޟ����fj�P���Qj�נ�&M���X�����j��	�<�wK���9���<�I��d���������t��%�<�x��Y٪�����h���f���_��x �jB>�:�m��.QI�]�������<)m,���M�����Q�(��(�s(���nN�HL� �w*G�N���PIf���ߒ/Eʉ<ϼ89�s4l/ī��t�W��ҿ��9�����X|�����W&|�cFZs��.��Ħ�N¼Ţ�"�'�H�>쥕�M�Ga���l�r��[.H��B��y.�)�������nPڳ�����
|��� N\��L��k�����|��Iz���֬���AUj߇&���[ I	=���3tT�v@9��$(8��L��HYsA^�i�fhsyh͘�0�*�f��S����y��U��^���}���A�KR�u�%�{uʻ��{C�G�B�'j'.��)z��3J�i������y�Ѿ"Ng)�p��K.T�"N��&��X���A��.�����}�:��NwLwD`i�^����ۯ�}�{�V�X�%_�"�c�9+(#��=#�Q4�� ��ˇ@�	���:]�&�f�j���I��
��H�Qy)4��0�1(��3��Ƨ�C-K�Ɔ��S�����#�'�^b���t�Th"]Q�u3����Go�a4dPI�"�|�k�h��5I��~���|��Mhl�A;OE�CV/��8�'�X�2�
۰�"f��~%2"}k8���7�ؾ
��w��dJo�L��G���DF�p��j�u�7�r{�=�J���w;���������X�(�S�&�a�k��F�����J��l�'�����O�Rp��Յ`�Μ�61�Owk�scdD*#�9�Kc+T���[/!+o�ź�W"D��������/�������0Ԃ�����Q�] �b�b����CO�3G��=k���@Z¸>s2)@�F,)	�L�:���� oK�c��*rV�o�${yy�KY(����9�]犘;Н)��/g�:RL�ȝ�ӱS��=���О��6���ux7���P_]>ې��)���=���{6(��z ϷjW#�w�6�+��s{�ln�km�QM,���my2|�\4y���R�'L��w(� GH�N���v3�-d7}�J�i��pᖕ�x�a��9pP�����v.]�����4�3���;�m���~9ֱvWb]�$������~M�z?� ����CR�kRhY���C�jR��nuzX<P3��8w(swC-�fz�:�I!a�9<]i>tJ�zQT\�B��>���0z��n�j*�k��\p de�H��4K��L� �]�q�t�b+q��?Q	)��ƕ'Tps
�DﺈA��SD�\BT_p�6� 1�i.@:A7��>0]Q�yl����m�h�l�!O��@��c^"(-�]�檡�YNʲ�����㻬�#+`s��u�(��U+�b�
�*��X��h>�n�Ⱦ�&����Klt��6E��ٷ[U�.�rb�䲆:��|M���%8�\f�����k`����<�V��n��Sf��\��k-j�~��^��#����b�;&��a-�NJ����,I����K��2DV(��0���+��1���D�G�|4/#nky�ԗP-x��vy����(��LOW�Y�59#��&�X���(�G��*��7�|^C�sє�֐_�9ǳYP��"���6�~�xI;޴�ɴ��aɝ�uhs��y�r�8���ۮ?�t�)�/,�!O���7߸pM[y,��,������dW\9@6��Sj�YI1�3��
`v���&ȯ+�&�F�pA�0��_䠀���P�����Oe#膘u���W ����7!j�|��y�%)�;���}��e�C]t���}n?��H�4:�â��9aq��s#d���@H_6�J�q7A�bvV��)�Y���S(a�������HwE��T�xa��s�q��;��U��!H%N��<>��߸�ZϢzt�{4V�5e�;��r�Xlv����@��k]J�9�SΤ��ԛ�W0����@��S$TF픥���%� P��r�R�=� ;L�W�h$���S�ʶ�!	d^��o;3b;��383��Ɩ+���xBVٙb���.���D�"�w��͛������@\Q�a�8p̀�
[��m��k�#�ے'�ov���<�Mp��b������>S���uء�Z��꓉W�j�R<��{�H���o��wt<�V�j��Is�f���k�mW�BQ>j:�n!b��H��ͽo��m���"vR\�c6b��A��Ԉ�[��vՔҗH��e3�d7����7)��}h���Ơ��m#Z��H"w�%o��j��/QLa���|��o���ð�V��"|/M��+A�\U��&k��$7�#���C�I�|�͝�g���(�@iNTr�.>�@w\uwn��1�(�H�ʜ�͔��}~����Zz�AhW��Ȳ�vQ�\ �s���@<�����dg�����×"H�؃30xq7��=�?D�������Z��b�i��=|ZO3e�����o=0��>�P���\��yG_k�ز�n�s�
��hΐ� zw��j�����۫g�IW��ɱR���xx�*�_gWJ�B/A"����8؄��a��ݛ*N?�6���kC(}P��cpNS�`�߸aΆ���S%]�1��?��hV�t-��"���x؆B��v�՜1SS�+��-J���\�(�S
m7����N$�����o�F��^�]�t�~u��JCY�˩�ca�i��g&�,[�(4K����<���A��61�������E��g�
�]#�IC����>���-�Ur�nݯx~o2z>�)��afH ����{�o�O3 �^��ہ&/0���R����0�>�گ*��_�W��{��>��л�X��Ǻ�AD���M�	Ԋ��I���Ou�vF��R��E�E���Qd��c�a�P�ʔ����"�M"j�Aܴ��Z x>T�2T�F�>�>��f?��j�
��י,���({s�td����9������v�����L��{�}~fwr@�����裌��Tf��7�+C�֗6�\�	cV�`���R�H?f��V2�x��m��pY�H�LQ|?wڢ+�L��=�YTKbc����0��L^�����rީ8�j{y�S�rw���
�����8S?}�~P��,Ex/C��h�kg��k������8R����Wm1���x���Qg$`X�8'X��=>�t�?b��\1���݇���%�Cx:n$���Ж!�
���b�@B�}1x}c0�Q��a�{���I�&{2A'�+ӽ�pw(�܇D, x�,P�/�_w�2eG5�mU��8�_�4�i����ݵ�\�}ZP>���^PQ΅(M�Cf�z;�.��Sfw\�IO���γX�/*b��.�]���Ƙ������������l��a�7���PFm(㸎ĈHd�������U�4�ܪ'�`�Yq;E�P��D�@�)!�f�@� b��D:[�⅍�u;��w�ѹܣ즒@ݍ�l��e��p��xE����q��	�����}G[o���2w8��-(*c�ӫ�жUj� �>7�l�R��������g
�,L?���1àdB9cN���e�������\ק�+��F��i���Qт|�^�sQ@�2�N�[\��UO�^o����{�Ņ�a� �f�zO��2yo����?�WF��欯['�`XM��w���{Y�iCm;8��o���<�x��i&������4�Jo09�4�y���A���5%�P���4Ǭ|y�,S�X�z�կ�!�$���ǖ�p^5!����O��;Ah��"�s+�A:��U���:�Aii�D�͇i�Z�R�-�h��q;#.����}�ʅ��_���-�sto�8 ��~E�����t�1�kd&�F̩Db��ȇ��7-L�O(ۅ�g�q��#B��w;�Չɨ�h�����K?C��#��%szL��_I	_��6O��}�\�m�<SUy|h7Zn瀮�������/�+�6�t?�>�`U����B_w���ZZgQ�m)�/�]޽��%�h�S�Gy�R�B�;���H��U#�*�ѳ��\��r��d�����o��l._C���8��BO�m'a������,�3{&���Ι��Ϡ}p�m�[A35H���cg�g��oc��v�sl�)s4c������ T�:3��ה�����NM'h�A<�(�4�aX���������zOv&�WZp�'Vi?�P��e��63'���-��[�����?�k��nQ������_G��r`�PT��9]�\�0��tK!����TrI8QT%��.ґK���{�WS�4]y��Q&�K� ��n��zn���i��j� ���P`��+�����4�݋�,-�qGK_p�ա���BZ-�j���8�Je����6�d�	�;��h�z���(Ñk����2�a_'q���pQ�~�L���Bk �Ƃ21�3��A�]7G��|�V�TC�`ڰW0�X�ܻ5`n��#p�*�col�-Dd!�N�����>/&���`�f�!�M��Y�Q�K��=g��e{�h�4�Q�����>\&;޷���qS��F�b��!�Pci��	Ͱo᠚d���fe�&�<�"�qӉQ�<Heg�]+�!����m�ɨB�@�����;}pQDS�h
l]��lh	?ñTl��U93��:�֪�ZXݫ��y�K\A�%kbĠ�pɿ﭅�W~p�պ �LIkƂe�4�\��$�ɽ̧�·>���b�i�Ց�k%F����v(�_ ���
�� ����`6e�h2"S�	���Q�D^n"��^��pyBSy%���oܫA�Q���!S��\� b:8}W���D�w�dz���&M��K�ب����Ƅ��!l�+t7��RQ���,NϧW�=bs����,[ <���4�0����R9��#V��ż�d}gU)tz�֢��Ӆ�=Ůj||����
��u-S#2�-�C�A�YV�	A[q�-��.f�P%V+/>Fo�#�Y���c<�U��#a:y�����Q�)��0MQ��'h�ѷ��8EG�IU��d�!7Z�X��ufE��6:��d�a{�:������W��z�� K0|�ʴ`�0��/�^��J��#T��3qd�xb�e�Y�O�`7h~�������$��r2�mb�x��JZn�v�(>;�L��e�֫�*���OM�Eҙ�}��t^�?�B�)*���m���՟;!4I�1�71{GO=���J���mJ����5��vp�X1m���vJ��퉅�c#���#��/��G�͡b��:a�RZ�%%I2{Dޫ�b�T�|��D<, �%�i9�VW2ˉ�f���Z��ӥqL��6|(�4]�N��X�=�«�.Ȏ �h��I[�waGs�z�\�J����Ć�L������\ˬDz�+FT=�P\�)r�p��uF̢f	���k����X�7i ���JvP�KmL9pׄ\�~�ڇ� �E���r*��(����X�]O���fg=ܘ���P�B�X�B���H�E_����G�:�w�"�${,0t�0�����ۓ%�|09v3�'�ɐs7X��Qڈ�d^%��sC�� ��J��`o�Q%P�)�� !�{��G�4��t\�7}/x����C�A��:�ʡ#�.-!����^��t��#�
�$��z��!]�܌⒜Ϣf�XT56=��
��]�]�M�dG�l"�1�_=Y��
�?��b�AL��W��cc7�į9�˔`�x�ݧՀ�X����O~`Qq��s�v�9��~��1i1�N�P;ϩ�P�S��>��L�	�i:`�����ٜ���I���n S�j)�J,��U�3Ů�!�&y�t
���j5�@_D��b��r~�0^�.zc4�af�P�����O\��,B� ��-��)��0�3G��!���M�3�cu�>��0߅S�n<�Xzge�LF�O�`c4���l��rwyi �۾B���mLIL<��*7v=�����S��eQ
ѯ�f�'�tK�q�]�#Nܳ�[;�Tj�+�\��EG�����?�M��O�-���$�T^�o�eR�
Ȏ�[x�l���e��n��%�=���ָBcN]ݏB��~Df��>�Ql�3$�c�C"�+�<�;�K��Ωf��)�C)7���!����pq�IAA�I���{Y�лQ�����ObR�^��z�_z5`���+�M='��뗁�v�����,�g%T����������U�̳�F���j�B��u2���h��Wy'�$��_39���=:�A8O R�&��$ǡ����*�gs���߷�T*Dn�Q��Zv�6C��/G�@8�����Dm�_����Xu��i��l�1�����'PU4��U����%%t�<���Z���C/�1S��<M��]�$�@TM��e��,>�J���vxpu��8�S�q��C��CJ!CH���X�m�2�Hg�1�E�Eڝ���W�� �闑�<]�M�F.�΃7�2�,(���W�l�ҿK���hG��`�;�n'9�A5%$��e���HH�~ T��@�Y;g����	��NK/~2�{;GA"�k�Ɵ'��}�yT�q��b����6A�儖l��Z5�t�����<b���h
�_�&w�₣"0x�qH5 ȱf�BO;_�%P�V/��%���&�U6b�t�� "jr1]��Ш�a�6�f� `Ww���n�("�k���#@m��/%.�qęi�����$��osC�@msUf��|;�Z#�ea0��`�gS��"�H�/�)�iL]��8j�t#�\����U��m� 8fh���i�ۢ]�U��!�n���2e'�Ok��]�sif鋗@@���j=�-�Jz����ê�s�[��;6���΄5�\�?.���T� \�oϲ]�=���]5�b���������5�[���~~SƨY�����H���.���a���k����ڽ�y�m��� �Vm*|!ףk����3�����Dg請�yF"��}��Q�/`/E-��COb��FArS�J��i5}7B��1��kZC���hc�Rs�U�<^Nm�LǦ���_����g��\�av�h�.�����񕰳$�KF!!�A��?&\���ia���?�-T�t̍���#��'X[��d�L�Dk3y�.�����8˽��NЌB>砸Ce|���A�x�l�����r�E �{�+Ľr�bئ�PMC6��n���׺��d��cyC$��74��0P�
�-����:�*)4�Ҹ�Y�����<��Qj����ՅxIbm��(��l'�^�+z�M/u�2��i,)i)2�t>��[��i&�$�'�_��u2rE���������l�� ��8]7w���(Jږ�r����$4U���+FTK ��#�VO�����@VN3Ц��]t�G��}0I�=w:'��m�.���@�<z�Y=y���9=��Z�d�Fu����!��i�s;�~L{%2�##W��d�򐙝g���X�K��X��ಘ�"�9Y�����r��i�x���:��1��yÓE�������#f�Hl<�8I�a�?R����R�怚#��]������Ǌ0�w*��� �h��$c<l�!=a�Jn:�Y�����w4v0��ߒ�j˅9Dcw��#D���s�nc�S�,���jdU��f�Jۜ�\[�뀢��� �XLi���~�%%��v�؎��r�� �@��z�g�{vIYǝ���2�R�L*���b�Y����;A��T�f��>��s�r�r~Z� �YSĔ69R*5�)T����{2{��9��7��`��4(Hz��2�pL��r\�740W0W4Q��^��Cp���/�1YLEU���3�b �}ok�d�X�U���6Q�_EH#�sE���g~���Z�,�ّ�ad��[L�5�9.�D�xj\��7+6lJ�ä��E5]�ܼ�^���޳��\H%�����TEO�{�E&���o�G|*1�9m��&Y�?��\P�n���m?2��Ȝ�����m,�4E��͔���.UO�Uș}��i��G�_4V܀�af=H��[�|)���D�?F�u+j{)ˎyhw��g�U����,_�)�rl�Y��H5�
��,���A���5gS3UQ_|b;�6���S��t�QTZ�
F��ƈ�dގ�n<_Kl8��-7�|�����w�3�&&�����2/�� 8I�t�]�(LIz���c��Ci ����&-D�k	���x�f��F��NmlO���ҿކ͐�\)�>)�ǝ0�)M����|۪9��'�*�M�2g��ł�@��|�*49�}�'��Cq���ڟ��@)���?c!C�>��,ՠ� ZI�]��v]�L�И({u�>+#��$_�^�;0o�-}0�k��ab'�*�@kMc�m2�� ����b߫��1��ܕ�C�t��t���*�%��64�~�>�_/�c��G��Nj��� �/zu�e��?��!k ̞V�������z(i0?��'7m=��3���:3%dE^esDaH���K��CF�X�`���ܧ|]��V�I����Ilz���?}�UܘJwXΡx���ʩ�4��D9��pa-��X�!��[��u���iDˡ٣$�-��?��I�(̷��
�W��� '�����oO�p	2�8�ň�U��s�;�٦_����f@����~�P���cD���6�,��ǡ�< �_K5�������&|"������~�&(�(�
L}�P%*�B<Ԫ������J�w)Y�I�ķ���