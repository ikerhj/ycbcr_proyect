��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.yu�=�6(I0Ĵ��P�]�~��er�)�Kd
{С"�qi9������D�~�T���p����Y��C?��ڿ���XK�U"��^V�I Y�lk+(�ˍ������6��vsx[
��3�$���$���������]��?35���3�Ö?�16:�=�_���m�C8��+��dN�n1:�"Z���K���Y��	]s���ئ�eS��讑�MN�����3[.g�rz��?P����
{�!���>�B�=��Űe
~UtL�������cGK$i��0BK��Z��"1W��¹my,|*/���}�)arx�]¦y�T[���oۘJ�(2�Os��"Q���@����b
|��ӂ�AO,dH��K�|_�lHL\2���RN��M����z�bM�}d�NO�T����B��Q���W��S0�*��9�-�<�����p2Lɧ�cO.!���P.zmZ��Lf8�쩡���!| ����Һ�b��P���� K�H�$1��F]�;�%�8��1;�3�>�sV'�:������MX�f㳳�I�[	�4�Gi*��"h����n��&9o�7��NAAW_gY���N��O$���Rj���6�u1��J����]�J��xOkX��b t��&M��@=��,H-��6�meS��>�ˈ9X�2��4���;D/�t���ml�v�l8s0�&U~A�*85�A~�[�MfL���*�<|��~OPC���#9]�W��y*�k�$�A��FK�_}�r_�������{���i�9�U[!�력������@�Ɨ
���p��u�`���1�Y��,֛����I��(7��?B�`jy v2r����&��W}	Ӹ�H�:RT�(�d� W-�9�%�O��KV!:�+�0�Ԭi3��1ݶ^bj2u��Q�J�=���>��vP�.k�)��eh
؏�G��l%����E�an�Lu�"�5Oa�h�S��l�����WD�'�!����;�l�����Q�gg{��8?}u��u[߸�_�-|����������J+X-�n��U�S|�a�P�p��r��S�1{�$Gv��T]˿��v�)�m��׋ �;��l 	��W�f ��}C�}Ծ͝C�D�Tݴ/j���?���v�ю������{�/�灻h������@(���Ŝ������Ci\���u�	7���]��'���JQ9�p�{�h��܍���Y�[B���9����eK�u0�c��(��4�x��1��۬��r�x?_$@�)���&G�%�@֋�TY����72��sʇ*>��X}M�r��FZ�L�����M���Zw�� ��JX"qv�1����j�[rA�ܡ��5z�/�Sjh��������T�o�h��x^��8,�i;��
�(&#u^�ɳ��4��d:�;��\�-i���};����7�n[k��3�i�Z�<E�¼��Ef�%8��5������|_���{C���G1���-�y���r�I]��p�	�+����Kꊱ]���в['�N�a"�bN,�o���e�l���h}6*V�Y���2���}�v�zN����ܥ Q��~���Мq�lt	�D�QX�,j�Oj1���X���CK�:p��-��������m|��J�I#� 3Kd�`]Տ��S�7�@�O	��y������K�b-��:Pp�hFcs�c����Yc��i�Q��\��}��[;���څ+�מ��inLTd#'>���8��E]�������$0x�#H8SAD�*u�r�Q��gF�z0��;��ǡF��:�C�;�^9�#Nmք�Z�@��b�H�?E`l.m�<�����6 ��uA~�1�iY��e�����Tm�GR/�a�v�P�|U��z�\'�����!=�����$2">7:��4T���\�c~�����]ݼN�8��� ��qkc���P���n��z�")Z���
��%�}�P�J:�)�W�������H��#�S�D7$��v.�{2*�,�OLG������I=���ke�jJ��^�h&��vƵ���4T���z��Q���a~��.S�嵦���p�?\O}�S�	x�����é�H�W6��Z����
��R�2��F$�2��E�N�}@�{�@���}/X� ��j��,���~��'�?8B+�O��U�ղ������.i�j�g*�;�&E(���Y$�����&U˽!�qw�&�W ��}�k43�^\�����ڃv�B#U(��M����X���D߁��8����D��M���#�I_�����c��	ϚO��c�D|�Ҍ�����B��M�,��tb��0N&�r�3λ2�&ѐ�[u��T�s~�
	�$*o�QB�����2g�XV[�;}ݪ�,��V�/Z���!�l��%(�lM�YI�,��{��ѩ��f�/&�sRz�S�ї�\�H�E`#��L�8���v�S���_����5����%,�@p�V�%��3����0S\�I}��=-��'��!�O�. ��#��6�2��zt�^��)d�]=@=1e�|S"���2�)�����K��c�An\r`9J=��ҟxN}%�Ě�y-
~܏�ǜ����KKeJ}7y�J� �^~,��$�f��'��VF������H�%^H�݀"�BDr9i�IataЉ�g�8)��!]�3ym�'J*�Yft�1�E٦���!<F��QRc�U��*Ůc������<��Co��A���B�Z��.L�����݉�<ظ��5yL�a3�2�6���	��p��>�)y��26��)�����]��0?�����qq�:셷���-�1��bR�$(�'pޣ�r��B�j.r\f�[����S�(8�R���i�t�N�N���R^@�r��OB@���wsR_�T�ӊ~�.^-�_"������ �&�x=�}`+j	7���[�1|�C�o�2�����NW9�!�V0* ם��&?�2� ;��|J�~�� ����C;����w�ռ���D��i�#�=|��;.q�6�7�at8���5MԾ��l�Dw���S���U�J0H U��?�lt[����!3�H�Y���%��{0@��V�ՙ�z����
ZϠ�e��,ڳ����o���1q�� X��&�O���AG[+�u���$yڿv�	��f^ '��Ҋ��V(hP�HJ�/Sǯ���R���^�V��m��M�y�[�
i.�;(?Ĝ\�	=�XS�Z��a�l��!.w0Y�[�}�`B�|0���@�x��<�s�۷X-�-e�= �-B�I���Galc�֯8��`:b�n�8�d$f���U�E��(����ض���n�7�-���X|�x-*AU�7����@L��:_�'�>� �F��A�Q���W.��~��Ԋ��]V��i������8w�YD*��W�e��-�@�ʳQz�ɪI�+jhk�QM���?�����R��s���"����U����	��I�؍i�{*t���Me}���:��K$�Y��m�tn9����]ZQ�D��x��ݓ��o=�: �0ҶWqA�3��vĎ�Q�����5�Ѣ�˩w�ɞ$<$B3(��7��V��8���
ޠ	�|Vz�h����~��қH�s �Z��Fa���q���y�����q�q\B�49���=���li�SI��F�Х���`)��=�����ђ�0r]3�3[tZ�BN�࿶�L�"溺�Y O詣L=���j9����giBt���k�W��j�O.$aLx�sm!�2�V #�1xt�G���H_���	��ǵ�ƿ.�q9��1)��.�<J㢡�?��jk��{=��\�:?�6�*Ց�m���������#�6�ǅ����wP��Uϗӄ8��0��0����{�J`ִ�ϥI`�#����t�U�k%L��R.�vuk��]�x8�&A�(5��?cJ��B����(���D�HY�ޥ]T��`S7����Ufa�.�!��a�=jxwe���~����A����&��|39���ss�A�ߥ������i���Y�S��`�I�f|���� �VD7-�uG�Nʱ�/s��^�+<����*]Ջ��)�|e�0���S�7�i�����1��i�>ugD��S��e&2pExB<8���g �Q[=|&퇓�J߲V:��!7(TQvD�X<`��<�ˢ�����:�z�Z�{�z�≘�����D"sXA=h��T�:P�exd^��D@h�j>�N���v��J����~�W"-�_?�����>Z�:z"����}�e�ȅ�x��8��dW�C��և� �ըW���,�k)��,����� $��,�R=�i$�A����*?���5�<��+r	X2{��x��S��j�g�J�g���^sB�E7Z1s�U�}�&��z@�s���[+-�>й0�?�/�:ӧĨ�0ޛYZ7��iX��jur����nk�J�K�<Z�u���qu&&����<���s6࿂eZ|<	N�E�֟3|�����wC����,Y����ǹ��ƅ�&7^����x�_�G�j_�R�+*�]�G�2���v�K=M�hD��B��;K�f�^�K'�o�SB\�����.���$X���.�?Ԥ@@���ܞ��>�;�F���f
t�]?Z������,a9�^b�/��Vx95�f�&Q VT��M���A��%�P	h�d����rH�u�96�t���;/����,`���ME�B�Kw9�Q<XL���
��X@lܶ G��Pʜ���ӷ��hN�[�an6�˒v]9H����C��h���r�
��Q�ŀy��֓^p�b�cʹ�M1#6*����#�	�z�>+��(���}�m�[�T�������G
źz��"�QW�T�a"�Po.�!��-��_7��1���<�XL�o�e��|��ݫ��h��@D����k5g�<b�һ͉���TA!tfֳ|v0��T[.+u�o�S�:���v��J��hԋ�G4M�#��?��/��f��u�����mW�ѷ�GL��lI�����8,п1�m����Gm��B������Kc��e��X-�b?�y [bqo��co�M��͈P�K/�']�f��wVə���e���˼��X�*p�Y��|5�a��i��X��=6T��wRO�,~�|`�;�6�����'�,��f��(��,bE�v�I�;Ԡ�y��DuF7LDY�8A��-�%LYl���[���� )�y6s�Ɩ����r��~��� ���R�r���(��x�������=��#�RM�'~@��
�vS�.t�.ѯĥ��A��Z����	R~�LU#?�Z�ں���;q�������b(uu�)4�J+C�����V#/�SdF
Ǡ��B%_R}�m���;sy!��,�[z$�/L?+`D�̚�=3P�jn�jۄrF�w��\P<KӳygTb���*M,����;�؟��P���Ix�ut_�~1xR��u;FAO//G��7I����ܲT�"���{a�q�u�[�]*�b~�-�T#���sj8yiu�h��֝k珡|xMi���m5F����B���`n�\�s;����ܡKo��À.�dA���*���ҸO��e�]=��E�>��,X4w_a=�G��äes�j���\@\�h��'���"��+G�)J�&��a�ڼ���^����$�#Ѐ���B�d8I��ذFs�r)*�����1���������R��E謁�����1�Q/��[* �`�᷐'��ܴ�ˮC�L�, ��\R���7�F��q����b�Q�J�r��}� y�)Q`�ysF�\��.�/�T��0��G�קQY@�h�z	`our�p�u{�.�T2f�~3�S{T^h���Ծ[8В��DB���h�Q��э̘��,=c�u��fM�ޖ�)�zJ�u'׾ʫ-yc�iZV[��>�)����r�?e�y��1!o�-���8�Gy�!I_���z`�m`����?�
u�V9�^p���ebۜ�˩�-|� D���.��N�zV�W���c��btz ��]��wC3P ��2RO�q��IVO�&���"]	9@�y�����8о�'|������{|�p5��b��L���BsD�����jj�Ks>V��}=}Z��%�PV� ��qu$������j�U�0f��dD�4m�5nЊ>�B�	Y�7��01��n�E�Bs��w��Kߗ�oH��}�p��MEgHf�U1���?�_�/~[_�M���yim�]���f60�.��2l?*����7�b"e����_�6
V4 ��ȧ���(��@�s����/<�����k����b�Q�˗��zs�5��Z��|}�X���QpǷU����n�c8��!��i!��zYݰ�X��SÉ9�z� ��4���Xp���J\�Ź�Q�S��3�rqd��]�c^%�x-��V���r^�N�zo����mR�V%#�&v�x)��cr&�S�Z��Y͇�!�#�q�Y�7�RҚ���p�BA�ҩV�{:B(��X\['���*���D���8yp�{���l�f2i���|0����,��Q���g�m����.����+B�n�����d��vo���)��x�풁��O:���m�rh�� ��h��D��N�u��D9�O=�����.~$+t��c�d����q���"Sc�\tL��� ]Z,�Xk<�9��>����٧g��?l6�_PA�M�ֽ��kW8�d2`�G^�%��،苹-n����G$��7�<c��OSjU�7Z`�VW�%�K��o	�[��y��Nu�#V����&gO�W�9�e����{��z;�ڈa3�R������0��n� γ��ѥ�W��r;����<گ@���ћ�5���wDt��gz�LQ���Z�\�|�=��`�DOy����5>�e�p�(��vK�%ѐ��U��y��TR���Kƅ�~Yg���V�U�A�Rd^�U	��[?��EBVR���Yf�Rd��Z\�w����/MZ^����N5k)�޲	�����W��V���rP`HHKh�P�<�
4���(�#��Z��QhD�r����ϵ�;�n�i}OHfn��#���yu0;e�qM���3}���r#[���n=��x(�,�lY��)�	��
9ZZ��S��=r�>�Jie�@��F�C;]<�*��<�������RX�:AH�s�;~����7�c�-RԵ]�����7�X`vҩG٪ܼ*�����~���$;%����未�P�!��W�页���c������
�	��nK7�5�%.�� �+f�{�y�q�4�R�<:�?�Z�l|�j.[#Py��zݪ^3�To�B�i�h�xuD�V���:Ќn�Ȏb�_Rl�{��A���ȳ�!�!�C�oa�m�m�Q�q���E=j"�Q�
���KX69�%E{nb�º3�ض���-
){�W$%
s��GS����_��A�-_$Y��]��zM��'��D���c'��Nu�6����'cq�Ҙ���F���6��#���������?+"#!��ϲmeܰ��لPJ-%*e�[� 4���bّ�@��Ҋ��h�D��{&M���Bũ��"�.�gZ2��yF̩�9��d���#4�5E)�_�Ru+C��w��������ףG!��_�M��A���U�٠s�뿝KQ=�g)!S�[�fk�\�XG�\_Q.n�"*�+��oC�V�07ю]:��ۙн�5��x��Eaʧ
I���c�eټ��g�rp�F�Eޝ�5ȃ���x��!�����L���!>6���S��Z���K<߉�H%�/���	�b�<̓�+\������ԫ�<���]\�+�Z�y�߷Z"�Qo>�t|Lj��"��G�W��b>j��Tp�w�-�Qi6�@���b|nI��(��s,ޑ'���R;�N��D��T��B��#��+�?4H���AH$.C�̓Ն(�ǜ6��VZ��I�z�G0)��YR�8�0�"ť�m�8)5h��o]�S-Ϭ����EZR& E��O���M��?$,W��\�
�޻��?��̏=�!�\ěGd��v�Sas!�:�x\��z��J��!e
�x��`Ҕ��'o��q�6�d��?zx5�����Y�gf��01���-�(���8�0n�>�r��$4>�D��� l^�R\1�Je�4���'�������:�f�Ś�5T�6z�"w)�����Q:�fP?W�[Gk|�c� )��+�i�IF���d�\{u���c

�&����7��Ԁ"Q�pܢ@���T��oKx��4��h��p����,L5��|��D��a�p
.�/u���	b�	�����1��8x �I��x�RǶ_�1U�G��pN���Ӏ{�q�Ȫ� x��r::5���V�)�ӓ�vCm���1����,@��S1�|�_�^��%�/JF	�#=[:��6;{��q�b���6�I��9��D���	J�8˓]��B�Y�=<x��i��U��D?���F\o��-�όR�S���^6�(y����#�d������z9��%ƪ����+�(�=ŀ���4����HL���͈�^��@��T�E_R�uG�:��R�F�yV�>��;�K����Q�I���jm\��)ϲYg
����~�F�J��ic��oJ���Rs�BQ+,~��5s���I�w��F�J��
����_�Z����	�e,�ş���0�oM_�&��6氆sJ"Q�N��zC�v��@ׯ$(�VT�� ',V,"� �Ř�qKiU���8�v�g�.0h���`ۿ�����D٫�@�ȋǭ27�D����qf�6��2l��K�=v�΍0+QA��y�0���P����s�{ǚQ�С�G`G>��f���	���uv�gu��d׸��oDq0��9m�M�tr.W���Hn1�& �cNmr�l�b��asІV������Q�1��}䵿z:�]��v���,�;"��+F�#t�j$5�Tf��xږ�<�{����O,�K_K:�IZ̹�_��mR���s���I��_X��IM3�b�8҂�+����+���c���ؓ�y��oW񳱅��쑧G��Q'[�k��A�;$��[د�PPŒ ������S<��aJc_x��cp��Ng|�*���s��+�^ȘJ�������P�L�f�y�U&L!g���j]+(Iʍ���f�i#�$���G:5c�r���������ă��y$`1�d�A�=+�8x���āB���Uz#o>J��K�s���Y��&��W��bD��e���42�]Q��ϹPT\X�
~�A"�0Q��ʪ����)V�����2xE��w�C]jɝiF�@��z%~>��Kۺ���߆R6��� vs�J����b�9���s�V;�Z����q�w��O�!�#�I��r�L�-=�����|���m|��O�d~�o�O:�����43���t�7��;E��2�	,��k�ٸ`�X�u�͢�q(� �'�j������Yy �$�1b�x�yޗ�5������:��P�ˢT������20[����5Q6�:�R84o���	y�\�]�`)ON���%����n��LW����t���)���g��
N�y�C�����q�:_�\\>m[��=9H6	��6��V���み^H����4]L����14���~���àr���yj]���5	�g��{y�|�>�w)��i��������a՜�'vOn[�W��/���8��:���|ǫ����@ި��1����r�o��9-.���bγ�TLa�Bn��U�����T�D��6j�C����ĺ���i�V�C�G܉K��|E��0fuE8�c>D���܋,�߂{F@O�0p�� ���3[��^���O��Nb��3�ux�E٠Ԍ��I��c/��e	b�9�Ტ�N�3P�B�����WvR�]�;��7�xm��-��|&��1j�
��5n�Dޱ����b��+�_�q�\�qXX���E�
r5E��\�%�:�)�����gz����l	�L�.����s�����<oS:�u{>���cTA��J��ב���������o��ǅ��.��$�Ȓ��)�撡�<U�dL�_����hF�d����)Rbw�#�nȀ�a���,b�(�a[%m!�5"��G��$ҽL�#��@�#�M��a���/ܾ�E�i���,������t,.V.p���G~@�/��/D�,yp�.�)����z��էG�B-�7u{��P�3:��v�<m���_]Bo��
}/����C
�܈�Рa��Ow �Np`R?�6vzM��i��С~ei���Eb0ҩ��*b�!֗Y��������q��C�]j�z��JN̍y|�|R������e�=m	|�.LTG�d�%/�u*82�'��a� ���� (T���/�^��פ�����N��w�]�%�+��t<ӕ~ھ�3n^z1��o��Ie�/�B���J3(�3�SF)���hi�i`��q:�S|r87E� �t�Q�nP@U����uIl!���oVYU�'
�,KZf\�2V�|[��y\_b�A��T�!�3�7N�)�1/�]v_����Vm��f48fO���+��H����`�*<���e�5r��`�`���-P�yl�(s��o��?	&h;�Mϴ�R!�����I�i�Nh���c�۸ELC�O��&���r�Z����j�î_�9/�4l�|ɰ"���S|��`<���g��mÒ���sz� �Q��V�W�׭���꧎�䰜�5%H�1b�s���}~��h/�PЍ�	��?��2G��̥����|ӵ��*=�1��5���".�u�ͭ��� = ��\�%�|*��6�&.S���㲴q����A����Y-���I̘&f@���[_��P�0ivR��zg�����������q�P�Sn�7lu���֗�rm)�[b��$�] �1�s���Re��E{�]G�­��[��0Z�Ʋ|��3ճ�&���O���buD�� �
�k�JD2�H���"]��^�l�s��Hyn�!�ث�8f��s��i-��sP��d����f*�}����o�4vV�i ��e���=��?�:A_��O�̝TF2'u�m��7ê���2S������Xs���j6T˦�>U�#-�����~�P:�7������֮ �r5I�G�]���Xp[gZ:u�z����F\(8��pf~����ʲ�r�Oy��F�?��] ̒3 ��2���t�\���˳�14W�Yo��4��8��:S =� ����x��5�n*��3��� F�p*�M�-f���S���U��zR0��q�h!J)�N�����D�GJ�"��)o{�b��.��%�0���T|+���_L`2��!��Λ	�(���Ɔ�q���WaVXn�S�m�%C�cFD�Фko90gڄ��F��!�ݜs~B�b�r�HY�腁�����}ku�(��9����Y�[�!�-�g�6`��e��;�BB<0�T
>�k�lQ��qHu�Lq�%�7TY�hX
��d�4a��2���DdX$ߖ���$!X��~����*��ʚ���XF��&���� pj:��ܽR*m{ASa��b'�_�9�����e�_����n"i9TDr8�PB���]Dr���K�)Yw��dW��4!�%AK�daF���#t{����=��Q]�\0��?�KH^mk'���zB�A�♏�U�Fs�Oď|���������4�|xo��i�FMJ!Zb�.m��H?�'�(�^17�OMIV��f��jvd�P$ݸ��C��;�����ҝ�[$g8���əqb���3_\�/�Z�?L���8�WL�Yf�(�cG	�'�>��B`��-�l 9��t��m���?�Fn��Z��m5�}�%yi� 4*�P�V[^y��_�_���'��g����\K5`��lv���A�0Q<Ͻ���D��1t�������C���u�%o`/�x��ڀ<˺����..=��*5~Q���Y�D[V��I�n9T�<h�2���@�D�����p��ɖ�e�|1��LeU��W�uG�g�c��d2�!��aЌ}��
�+C
�T�,8�<����c9���X�{?/����uAx�+��+I1�f΍S�eII`�����w�>�����[g���x����s�����R�a^$��:O����s���-��R^�:��-F�\F��^�o4"m�_��RN!&c?�@�;P8\Ix]r:�F��C�o�rs�drJY�#D4��+�+��FD6�$&xe�����V���{�5EB�+��51u���/���h��L�ƻ>G�w���}N��`��W&���@]�St��U�_�1�1J\� �<�Ć5جR�+�f��w���Tϑ��'��{_��D<�>���O���5k]��WH���:�&Yk�ÃA����i����ރ=�z�aEi���iq�-`$�������e~1,���	����!Y���p-�"�*�szK<*�R%���ϗ����ٹ��Jm`���r>ẛc+�S+�,ٝ�fկ�8�v�Y���\o���2���/;�A6o�Yg2u(�!k��h�с(h���v��G�";G��������ދ%Yh�T0޳s�ҝ{Dw�)>W��4|5@[Ŧ_m���.zg�e��?nu=�ywyh���Le�bY�Ɋ\�!$��<>���}"�4�/Dm����l�����y�bx�V���4!T�2�5i����F]������#ęth���'	%��*n��:�{*��j�A.��B��!N�N�g�� ��I��|یɨ0'	i�v=N�������_u"9�yS�!�A�!,��Jw��/AA�5S*����^ɴܹ���2(����R�o]���T���#-��~yg�B����ػҗ~9�r�w2U��3��ω�Z�>�m�yQsp�ޗy�Z�x�U�7a1~���؂�*c������|�OX%�}��i�����A�O�˗`�D�h����N Q!��:;q���s���D������'1r�KJ`B
Q�yyt>���@��&���g�;�Q�c�^b���rߋR�FN�ٵ&���؞�謥P����z)V�����YX�fu�&{�-�ǫ�ܻe�}R�C����k�QU��A@ 7
�-sy؈�=�H~�=}�b,rxG�" ���x���:���=����Ѹ��J�ν<����h����uw��N����9nSƸ�p���K
ԇ+&�IZ#��M!��F]���Y��n��^�Gbs0pv�����������ے7>�v!�;7��#&��/�˴�͌0]��_!�~��h��9"��~�p>G�(�A�GG��&�W�~~��x%G�"rzI�k'�֘.�����˾S�W��R�O�d�Ї��lT>��k����9j���x}��+y���$NV�76���!�8��iǉl�<y�
��}�js�L�?��?4�Bҩ��I'�p��~��Ʀ���� �L��v�p|�< ߁$��cLq�u�Fs��{�%��^� &�9J`_���%���y�U�uBr��̇2}Cp����_i��1��	�k�ж÷��4Z�jȕ=H"E��M�>?X�{o>ʖ�?O�7�R-R��N���[���];�zH:)K����)�QSZ�E<���s�Z^�ƭHK�}��(V9W�tOϝ���r�.GX5H��i�Y����A���j�t��r-~4����6s�ӎ�S�hjxJÊ��K��ⴸ9cK��[	����r�r���P
���-��;��@��%h6T�"W���g�#�[+u ���xpSl��5[�H�-�O���Twݑ��	��	?�V����X�I�fFc�gX
�.�v���@6`(x��x����Č%B��U���I���n�=�
5	�KB4t��ʓj��s��7��S,�NQopl~R�j^)�e�V�+����,=�xv�Z�hi ������~Ne5���k��fH�҂�����	�9�+3���<ૠ�߼�-�/e�M#w�������;k�p'�j� ��r�rj�B��ʛս긨�b�������z��	y�)�D[/g
c[>�bi�糍�rQ�x4>U�=���u�%�1�o��C|u�|Ԛ�L>e=�]�����س�������+������]4���k�ɤ��]@eܡI����31b�Y����:4{�B�M��^m�@�i6e���Ј
9!K����YMo6mؼ�kÃTG�i��Q��*��	? T���P�Np�]�c����F�u���m�����:��o�+��F>�L"��{��J	�;5��2��i�����<_��7��\�kީ�'�"�B��-�A+t��F~ fGw��(y����eu|�Op����vw��K`9rP}I4���ga⹔Ax��*.�ҽ`��bӐ��J�# ���y��XQ�q|��6;�ƒ����*�@�t��������V�ȸ�j�.���)Ԯ�ch��9���ʣ��>��dp����s<�(�
������oA�jdub${R$'ED��go�%�@3~v�}҃;(��k�n�㯅/]>yg��k
W��A�\[����	�`U��.����, �������u4*�Ͱ���&�|��4����z��O�|O͍N�X`���8J9!��YdR�����k�c�%�k8���������{��\�?8�����s T��IO���� l��T&�i:��_<��������f��T�����),k�����l$��;��#�t^��?D;'{M�8Q��4���'�d���Ȅ���i��B�ߙ�y8`�e`��r���������"�G�8�$�Q����Z�ƈxla������բ`!V~��^��)g�D�d<8�/V���U��K3�1}��K��"�@*�A���ד�J��`^�D���4��"�g-�p���?I[��%����&�����3c�W2���4�!�#PT8k�}�L���I�|������:�0�P�#�Z3����"ca�No��Ƙ�+�{�
f�i�&`o��tP���'}�g�E�1���%��EB�ϗ�Jr�����]�E�ه�C�GӰ��׏=��\�4��DmY�2��@�Vx
x�g�x7��r,9�c�Uo3��4�)e}������r���\=]�[y���d��U�T�ͽq�!}��{��@q)��i�����BU��6p�A֕b�����l�0�Q{%\bOހaF����3"�?�eYko��AH�;��<Zb'����g G�V�AL�\�C�7���o��|���t��KqY��#�֛Ӈv��+_X����4�Z�(R������i�S��K�I��&!��ېT�}	iº�͂R}\_`�^��Ԙ��3/7��߱�@��X��~��KZ6���M��+8�#�+��gU�/�I�#S����q\j�B2�w��y�ȓ}��v�S�S5r;��v�?�]M��$��c�0RM5x���.J>�&��wO�[��~
�0�+y�H�-^IP���b]���ą܁k[1�|eRU�RۂF�1I��bg��VC3h=�+Պm���9��S6700+�n�6�ϥ�c��:��:2�Be=-3Wl:
���f��:Α��������4bɋ`s��_���5���Y�k'М<�� b0��f:>��D�;�y�D�Ȫ�H4�E`�9�t�.�2Z���y5F���pQM�C��4�)��2Ѭ��d�� !K�&Ș|
%�3�I�������t������8��`���,�X-P�t�q>on�`���%��oۦ��\k�xB����^����]�G�	��
�.�1)[�f�x��cDC�k,��U��&7�����4�dc���օ�>@Ί����=�N����8sBa{���Z{8%b���v�|��" � ��2\�����_=���	hc��jS��ipҶ��5��6�"dj��e�!S5x�ۦ����=���bZ������{����7��fp�54����9Z��Y.z<½>�"}2��t��#�I�2������[Q-z�:]�p�)� �B�H+1+��
�pt��_g��r�=��y������B����
��#ՋU٪�{��}s����Z�'(x�`8[�F#r�|���V�\���
�B|��(�X�oݭ��XȩW��U��f,6;���7
`�����K����ƴ]&<�������ǟ���ě���9 B��"�]�V�����P��p+_̵X|�Qײ���C	#M����:����y�Ԝa�!���'�@�{:53�a�K�#�w�xj�GQ�X����Q��Ze�X������'d���F��q/:U�GSEMC��EJD���֘�"��ڿ��dw�}�4�i���P��CD$�s�i�|�"h�ݓBa��.nx3��4�L=�X'흛�ڐ������M������=��s��Uq��)����P;���L"�)�ű^0���4���\x�bt�M�0�Y7O4�@�\0 V�y����$�?ۗXO�N��#{Z�b���=�?�4�ڥwM��LHP���[Ұ#Q�jf� �e�M[��όwu�
YxKU4���r��j���W�2�/΄��
�I�ޢ�O�H����.i�<�E�-ܔ��Tо� 8�	 �)�l��Ǝ�[� ���w�f�����LjG�K��7�1�F<L���eM��R��7H�a>4oҴ���%������H#�mO�9�U��
6qIM�p:jBh=C\��@d#|���t�������JS�^F^5Qm �P��dq1�5,ӬV�ĳα������'�h̬�	��&�*�Vv^�S�o>9Y+�{u���g�i��
��v>.�H
߈-/�[[��6�?�����r�݃ݢ�[Z,(���������B�n6mM�h;T�,s~�ç�	��d�$�_G��/�:�t����8> �_�j{�6�%qXI�`kH��i �Z{�[��u�iUn��NU�6ܺ�x��KI	���jN�󊓴�P��T(�V!B0�	PG����_c|�ʩ�mn?��L�4H�g�7���dE&ND�;�Z&�hm�Pu�\v���l�y��M@(���5ړ�ᓽk��en�Ȍ�Rg�G�j�nI4�ɛ��{f�̼������H�t!�E_bIVTH�S�c`����m+����P�C��g�U��?�&�ܾ��
�Z|8ބ�^^	/R����ӫ?�e_k�v��پ3�����U���g�d��xt��Y����ށs~������A;Y7���y�����C�:�+�8^�ј��ڗ{k�\��ʰ]��E$�L
J�ک�`F�aSu�f��1�,�̤�$�Gsi���7MM�OH�Yf~Y��,��dpK�6�|�?�5]���x�[�h���.e��SYm�_g�D[�8F8�=�\��c��h`�	��+i��m����2�=�3p�V{�E|�5���;���V�$9@�E��f[�:��hzR�JT���	6leS����䢩LNn��7
�ZZ{��N�}J�[�$*B	6(��n�N),&��ݬ�!��j"���u#�t8Gm=x���Gං���&�J~��MQU�ׄ,Qt�c��fb���3��qL�w��<�S�8���i� u���E+�;_�u3=>{�أ�7�ߑ��+����D�Ś�YS,L�#F\K��e(��&+VD��~�8m���	j�T��v��n�
��RZ��v}���^��T@f#����[�Υ��Z^W��8�Oټ��0l5�E}�R�����ihJ�)S�h)����L<�鎺�q���.�rA�x(=��9K<s�"��S�Ƀŵ�d��e������H8�Gbv�/�5��Y�s�F�P��H�CIěeʯ�D,�t�X}���٥�l�t��EegA�8�
RA�Փ{�EMB�&a��H6���h�B�Qy���!�\
�
c0�F1�JYCO�o�-��5��yoh�x�uծ�?Tǌ�������az�q���}{�R��/�d���,��%�����n7'�:8q���?�Ⱦ#�E���>��P���I�k�T�Q��gs~�P{�
��?RHv@��H5
�W��.����Fةq�%���L�
�#���!�����7��i)s��6�lm�?8+�`�4��$��K���&Ǜ5$2�@��­6�K��.��E�M�H���St�-�k����)!A��S�N%�1 �uO!h:�� 0Y�~�hQ���CA��+>mt�dʒ���J�N��w�����jd~^ZT-o�QEgѿF-�y����^�t�Or�=�id�%/rȅ��g_��Z�_� �m�w+���[�쮪'�顏�a�D�h�A���Y4��I���bs��g��f;��Sh�}0n�띆	�~�ܢ�#�#�$�͓(�D��pnw�W�!���_���k�a��pJ�H�օ���k�i��k�j�������z�f�%$�	�7qh�tF[{q�on����0�i�U��S�b��y����#\�?fӐ�.>o�=ݬ͋�`�I�|����4�z<[q������Q��:<�%�9V�-��ɒ���X���h�bk��AI�bS���7�I�=��$o:E��u�
�E��J�T�Y(�/�Ϻ���.����8��s@�9:"
���6��`Sb�2�تj���?�P�-q9���|vS6�y!���s[��C�W�a��7V4�[�v�|mY�jÜ8I<��?���g�'��Qu�`�a�a)�;^/�2�/=	Ɗ��NMѲ���PzN��$zG�xk� 0c��I�Gi�{��KS/3|#�q�*���ɐ��Y�?t�ăJ%4g� �����5����zX��ω,�s1^���Z4�h|�V�6,��Y��� �P<��v�j�Y̞X���-?�lm �@���N�Q4��Ur,���}�W�3��P�Z�Gb"�Q�:��捄��߆�'^�b#mb�(�;i-���id�#S�3_�����5�����i�S%��c9��':o���]�K��!jY{u������B���G�۸'���i�\x��@bO�l1��f��$�$�X�d���E>3���g�&���|]C9���m�\5V>�ꤻ�d!M��]}��N�� �z<��r7��V������]�������5��7�
(�B��H����(�&`)��9�B`���A�`Q0iy2�` ���b�襍�\p�8�Hu;��#u���·"��7���5hM��-燥!mt�d��i&�[�ZR�қ����Y�����'8�҅�S��+�U����dޣ��~�^'�3��Q�3m����[*t[T����osȒ�L�5v���[�>���1���ױ�PͲP�/<��-}��U ?�� �N�c��t(h��v�Mo%�y�l��P*?-3�Q[�vF�I�jm���&�LW)��j�:����+�M��7�W)�yzF�@�5w����r�tӐ�M�t׽6	�����~9��%_���y������<u�a�T�����X؏��b"Hؖ�8z=���_6.��F�k��r+I =/�����@n���m k���a�}�P��g͋��w��*�DU���w^8z������.X�D���:k\YT���LK't-c���i������H��%�	�9�����*%i6�4�駣A�o��`�q�V�
L0 �(.,�u���}Y���'!�@�m] ��_���I���"A�E��f��!�I%����v�;n˱��=([;��Br>!�6�A�b������B�l���6-��}R|e�F��a��
Z��1�,D�7G��0�����_�``�%� /���@�O���k�c�]|���)���@��v���BX����p2�ﯶ�=[v(C��Gȱ�S6��N�ڄ�uE��[+Ƭ-�^�8�T��ΫfE�i�>ٹ9[wl4>����du�`�fr�.>�D4fV.�
�-��Ԕ��/���=!G0V'f����KoDh7@���r��&��Ɔ����g��Ȩuw ZH�&�jV�@<qG�5���r�6�f,�gM�<�G+3ƒ�)�;Ӳ�A�X�EnU�x��^��uv�|8�Ӯخ�T�iJ�	�;}�>c&��!���k���W�D�&������n��~C�@t����� M�D�,>`|x���@c�jm��캱/���c�	��=�	N�58[�ex�������'}Pޘ%�J�Ux�&��/�4Su�*��?���=c�����v�p���x_V�-m�����������N�6���u�٦\+?�`���ϚTFF�K��J{�#x<Q#��������Oĺ�}8>��ѿ��n��z:O�����mD�|��?�\u�7�m!�r�WA�������dDUEJ�C�)#�>����q��?L0/��y�=W�W��C�~3>W��6�D!V��)�
��M���)�"Uw/�L�
�,�i�(��Snp��7�;4�'<�~2�OϞ�Ͼt�^(�I�g�bu���;C7��ĺ
��I+�t@�j�v�W�ɶ}\Q&��ߪo7H��͸���	�G�h�g�ub}U�S(��(�����;
�M*�3c��9M��d��l�۵ފU�~ 0SFWU��(|�=�[���kc�c�t��:'���qS@[����<�uJ?��,	Q\`@��=���>L��� p��Q+ٮ�~6� ),�����Z�ߘf����HV��l�*2�ƭF����h�/yw��/:��{�#��L���ةW���;��"��Cx~�&��]`Vw�8�[�x�5E,��e�O}\�9p:,&4Ѡ�r���# { G��eJ>�zB��?I���tG
��K�p�TW�^�F�2���BQQ��0&�-L3��� ���w�HLa�����l�oS� I���	��c|���}��ApWO�Y���*�ߤ
��ɤ��d�Jf[����V�+c���j"�����3%��x�a��iF�<@VD��bh�H���
R�j4���^�z��F0u�o[�Ѳ�&J�c@��0:��i��<�u�LjT�I��3��?�������r �����8j Ψ����M�U	O�2��C{�6�����`�3��.�<�%�QJ���K��R3��M��~IO��_������܇"��� ����i�#|���Uv��$�ѱM���Q�栀L_�P�d9��a��<��Y�Pl�-+] Т�
���>s2vJ"����~h$��ؼ��4q���6%���[�����lN�D�6R�l��'?��+v��qz��dYɯ=�0�����'���CV�Im�Q$^��~��տza��o��Gjg5�b��<|F�Y�g� �3u�uX�?��J�^Y��p�y�2J4�Z�=�1��S��g�ץz�E���������\�*���y_�I�	<�J�H��@�4�����@�Ka|����}�����UITm�Ԁ�]
�_@�g�ۊ�]q�5�lI_�@u�������~[�'��{u�	ԓ#�����n{�׾�j<&9鼆�rǠv�Q�ivH#��E�S�.0X ��@F|�85�J8@�\w�̠��n�� t��5�G�bE�>+\[Ew�տ�*_E���bY� �Z(��n->>�H3b9�?�����)
{o�Q��^�%\k9�r����VM0�fK��:������͙e�T�2��2���B{��כ����	Z��	����^:���!2t�����guc�L���d��k���M*�F ���U%��t��k��C�'1�S��6ɖ��7"č��d��w�=�|\1�(��r���A�//U��>� h��%4*�^��I�)5�ށ(h->�KoY����B��{a���:����A�x>3���q�K�L^oShT&�<D��k�ZKHB�/��q'c�X���#� j�,���:yA�x��kB���)27n0%1H���˥%]ڵ%E���i��P�4�F�?��2�	F�P�/�Wu`�/��#�ն�-V@j0��X���f�P*~�n0�g$��+���Tf�,��z���l?�㻃tq�2�YO�&�7�������6��dN47�5p�!���3�(���"�k�#˧����=�^�ceB�^�1���D�3Pt���m.����q�r�p��{u�'�c2���r�.��_笗�F*Rk�mS�zi��G[W���Lx�r%����U����Tٟ6�������2ZSY�aȢZG�m�5.
IN#��02�����W���>�3F�+��?0Ss�hn�z ��bNƐǈ���N���z �#3R0ե0�ıF�⏳ ���ǴN7��������G*�KP3jL	�#�4NK�(�T�@��'Pl���Ϭ������Rq$ �x�k�H"G�l�����B$��s�̭�e@:K�n.,�ܭ�<�o?%���dP<)��Zk�W�>Nyޓ)u;�t]4�O~6�r��6�V�CD�%��r�<y��D߼bi���ġ��p�~����2A�VtO�'�v���+i��$Ko��D���#��4"���/��
��N���g(����}�A��w��K\����/�4�3�q��s%���g9�9C�$�w ��3�V�ؗ�	��=-���0��Or+&���u�5�cm��c��W�d�Mm�;kDE��I�''ێ�����Al5��2�t�`[��x�E4��oF��a�C5��f�.~��ߪ"�;�>SWHLd��?@���E{�c���8 h��=򧄮_,ƌv��g��{gy�+Պ낞�?����R ���_6�]��'��	8�neJ��Ԕ�����?�Hí������(���B��/�G�֝M�͋
^^�J)��{��7��$�3�Ku\����p���\4��z���}���
K��R嵆�L��|��b�,Ma�����8H�l'�P��.`�n��E�
�La�`�����K��;[�zW��C�uUYp�����)��QO]�F�7���ҫ�>hEc��X �0&�,��BR�~�q�DJ_p��6nB�y$��R����ô����:��ќ٘�9�a�C�Bv'���藏á+�H��wG3u�8V4�G~^��s���(;�|w���5�ѽ}^����Au�z9Ca��� ����� �~*�U���d��[��?��z4%����
�J�Ąû�?Fф� ��:��jO�����oV���f��3�x�3�B�$�(^���z	�bwlbf�ג�ڒ���D�i�,w�/ww
�W��Z+��EU�%�ʑ7���B�yX8�x�V�C|�z�uN#+��q.F���`�DC��i;d�h/��P�Y ʌ��O�α:7���"��uo�yg��̟)�Х	f>x�z?{�4�,�d��)a�[����@7���k�4*��1#�&��)܇��J}���-��?LEq�����Ѭ �P��
3?讱C,{<�!��G��˽�ϩ�$o�	����ϕ�8c�����Ħs�̂�H�rw��,�n6����AI,���&����mlO;��=�f�#bCI�j���C.[�iv=Ӫ�����\�P��2�f�2aUU�گ�$��x�C�x��B�6��wU3��a��=�g�q���[�y޵�ػ<Y�s����
a��A��+t&� ̑⸹J�,CS�=��i�֐SC�G�\}�[�$G;�$1�'Tj��O_�0���sJZu[�.���t�7w�p���a�B|��l#����PV��T�/g��hF�U5;)KN; 	���_Sۆ��B;j�X�����r4��й��M��oo���~$[�+�q�n� �$PE�����H;/�aag<�L�#Ւ�:*B�C�-n����|�f�$ӓ
�7h;}�l�]r�ܔ@yL��L�#�|����uZ�k�,���o��!t�� �q�/��Y�>�h�_���G7��aO��E���i��%�p�Y�*�ۗ*�&q��\r��v	n�����鼨,�ض�F�x��2���[,."*��?�}����v7�w�?���	[�F��Xy�q�`
�r���՟ס�xD�R�΃�C��pO=9~�m�<_rȆTl7\q����r��o�{ol�/�,�Q��gI�uE�/�6-fF��N[́w(�����K��y�<�0�_�p����p��w���Wt���u�24��b;�3�Rʒ ѱ���x���_fܡ���wv"!;.Z��X�])r�o"H�QI��E��T���,����Jzn��e{Z���1������'��w>[���ź��<�z�n�T�g�&�Eh�O���\���'>�eNOi��!�<;J�I�N��@]�#b�~;�MG��Y%z�$��ي�y��er�O@岟7.�Q�,u��TV�`_���Q�ٵ�_��fK��b��eZ����<��Ϛ1�ATgw&&<R�E�M�P���Y�B���\�T���2��8�ch�	�E� ��dݢ��"�+�>U��R���V젞)�45]�|����x��P�pı"yQtwJP C)�,�<=������PB!�8�av����V�Wy7��� � ���>[D7�;4�e�>��0�.��Fp�u?ȭO�	��fp 'OcT�4�/�f/d5ۢw^�Z�-s��I���"۞%��0��3��p.�L�^�8�����~��)n�'����<��bF8z񭽄�2�*�
ߋ)�0�"t�P����J������Ә��(���#l�;w~�H�}{���Wb�JYQ~�t����T�3J[�v���M�M��=��m<g6Ru���Scѻ�!���ǐ]�ƛ��̗e���^�����IvK6HWr�*zg�^>��6���OF��)�L{�����j�_���Y�������qo!����� �1HÒ�h�\�.گ��4��i��:ɑ;�'y�_G���s�>5�b|Y,3���q�]�����)�Zd���I�e}�;DA�.Y�[�ssٯ��Ck�qk�JOK�\�b,�6��D�k��v��:�%���;�/��^���ͱ�䠞�����>uq9�	�:�;H��*?�����C�L0�{,���6^����1^3��"�:tNm'N�jz�}���~}|�\���9�CV�	 _X�<)	��.�9P��F��I��������1U�����w�&M/�a��I�T��bU��uY>E5U��*�k��Ά�!O��T��y�����6�ϫ-���$��\�3��tA&0��G
��T5��g����8D��kV��#��ٳ���m���}�����!�M��jzV�D�*QL-t�5ݺ=쓷_2�OԼ[ޤqi7?�P�x2��/ ) dr_Kz��q�j�g"V��<G���{xt�b$�b�np	�0�&fyG��>��"�{:.#�X�ױb��dS�sz��E�B0p����=�#�T�ߡEg�U��J9"��Pk�����A9ǁ��_���d��ۣ�R�E�_w���^#��-˼�,@���#>�o��Y_��2JE�bwhƼwA�/.v���т�-�W@dR�IE|Ա�Qj�w����l���οd��dz�x�������;���),����KI�� M���fy_}?�p 
1lr�-&O���r�	�1kN��*��іp2 ~���1$U������^#���`����A���ųwY�r��M`�Ww1/xK����\�=�����^ ����H���3����~��s�o_�N(~]��E=ոÆ����ݎ4��(�iF�h#������yN#=�~'Q�S���Vf��K���9V�N~q(�:�t+t̒K���^�)��)��8AQs<7� T6�}�:��=�}�hK��aq>�����t�h��4)�����zl�OA����ǀ/(C0�e�� �ڔJ��ަ(:���)�%�V��Z�W�k��L� �4�]�p-_C!g�\�딘��eR�I�����?���Z8�O�a�6	��z�"6��>��B�?���*ϤP�c�U=�lM={��\!�Z���!�g��Qf2���T?	� ��D�C�W�iD./2c��bxF�LLX���6������!�;W$+���tiw_��J��V�)�����PJ���IPc�O��9}�B�3�
�]lT��5P�zc�F*p�h>�[��/�!%y�p��?8U^�﹐�d1%V�p���0$�ή��/��7�X���@W	���u��ڸp�6��+R}��qD\L��kh�/ly���n�q&b\�W[��$��`�Ǫ��?��+W�}~�פ��y�/���@�.�nᑱ�w�ͺ�X��Ç�8���bC��Y��Q�����gg�γ(��y�F �9-�T��@�]��վ �W�F�mh>��H��H�b���>Е�Xj�R��<��R_&��5x�j�ļ�<���;1��W2�@�iQ`�p%�u���GqM�L�Z8ݵ-�!��h��6�=Ύ��-9�{�j�\?wo"�}#0M
ӲF�cql�f
�m�u�0�E���4����s���#g��vL�05U$��m�UW�;k�Ȇ~�?)/��G��I�\<�hD�|�]	~}��+��wg7'E_�0vA�jG�~�����\n3�w���!�o�؇�����@C�6�w���qF<)������͉���Ii�fUX�����jEP<�hf�}���!�a��j�P��"]J�������&�e��U��~4�s�ж͢�M��O���'������A�E�w��B(�ڟ{�X8� �	�I�K�ϯ�n����ރ4�FQ!L��k�֞9�Ԧ���"m��%9ٖj�'L%�a�2�I/G�����4tغxD0,��%K�g�
�
�t]�e�"�,�؜�D�16E'L=>�I�*u��w�&G�cͮdNn�r.2�ф�wN�i�����e���Pre�ӗz6y� 9MjK��qv�aCߌ�+��l��&~��x&�:x]C1_��~��?��[u"I��C�sV^�+tA�8&I�S�ǘJ�ƃ�g���*��[�r4FrT*�E?Pd���%)�9r�N,U~�/CPRh��UBX$�ʐ� D�~U��	�C!5�E�ŚwI#	�����Z�m;�<3XQ��us��Æ��k ;w�)��a	*��K��_��U�&y����6X��}y���_��d�bT�v�.,�o��C��R���*�������	�_ ז�4�[r��~>d�ۍ'�y�X��'3E��n�ߠH7��)��ڲ�L��}��R�%�Ͳ�@<��#��)�ׄ�V����[yd��mԍ+�{c�Ǹo>�j�����8�H3�q��| �� Rr�|bX������S�o�
Ν��]^zz�g�;;�C��j��'��g�F*.Z�
>=��3w	�۝��~��:-n����מ�٘fe�v(����R�h䍪V��˪`b%WOs�|�ȼ���B]kC�\�� ��q����(� �3�$��C��K@'���O���.� �ݙK�� 	������:���U��#&]��ڞo��~t��;��Q��'\5��e0?���st����K�P�	-ۦ�54����p��A��+�Ұ�� b�$ 4�j/I�q��N���|UI6G��rk"қI��"�Ck��K�g�Y�a~�Q�\.�Q\vor��+tX��&�,��4@a��R�$���?(XXM�E-�;��wxC��@����R���]ϳ��a��ڄg��}��l2/�q���H��Z/��lr4�ò�"r����=g�m�+D��/Gc��|$��X+���Sl�����+z�'��]��;JK��4��tZ�r�|�k#��^���1����b�Dh)n���c��t�����
=����Xؼ7r����Z6y\
��?�z�?/�7$�Zqa�-�鰒���u��(��e6��CX��5|4l���h��i%"�.O��u~)#���s��4oQ+H��u�)��~o/p�Oe��W+���wA��*��R?=�etlr�F��e���˩.Ի�jc��Q��o��G ����ʵ7�=�)~^g�ݦ�䃚�S��$W�u>}A���Xu�*�0_�j����I�_E�]��-"��	H�\Y���RS�#3(��Th2���҇�*B*d^�%I�&X�:~ �v������q���*M`����kMT�V/k&�'����A��ݬ�Ĝ����1����fp9� ��`�Q|�{[��K�EaY}(�����O��>��Ϗa�Y��(i���k/C�~�}˦}��?44�Rs�fʭ;�-��V�p�pQL�$��P�,S��V�f����viG��Y��2W�C����obt�:�̝���9���?s5�r�PPj �[f�����B��'�I:�w��1d��^�%�^/��js!wz�;z�����+��O��䄂�-$��y���y0��Cd�K�߄� n��ne\H��3�p �ˀ;��@��;����S.���fٌV����f���!A�j�0�|��6\�⭆w�TW�4��)�Ӏ��,�z�Y�ƻÙtG�9�w����z�vD�O��#�:�����3���ޒ8�r�&~��Fÿz(�m���}wqLJ�~Mm�$�;��jǲDdJyC��o���B+v~%������p�vhSe���U��Y5"}�]��ռ������m��@�|G�P�q?ޒ��y�&7��.	��ܸhǥj����p	�y0�ݦr�b�W�R�b(t\3������_��뀹j��ҥ�g���	�=���P����!Y��sJR�pʺ�>K���w���:]��5��0�"�_����ɳ��qNB��
�]W����Q��؎ f�q�M0�Z�o�6<Xw�[r蚥���&��.����I�jz�a,~w�7�]�h����1��s}J������eHЍ�)5�7�B��H?�S�e1��u�	�p���Z�ݓǇ�l�'������؇a�`c���@�2$}E���ͤ��9-P�\h$|��w� h�F��7�>X!:/�(�>����Ky�ivX���	�!���*�{>f��P�����D璦�N���G6��¦"��MX`����Qcw=�K��_P ����]b�V��;�ߕ�c��K��7 qt��5��}�6C%qJ6]��o[�Z,v�{������2	�J����[�͈��5��Rk?dsH�`�rɑ����w�@Kǆ߽�g ΅kb���o�I���L@Kԧ�8 �{ȖB��z-C����P\�ؚj�l��&]�=f�B ��=F�.�_K�lƫ�k(ر������4S�z��*�Ӻ���/��Ȣr���,�EAa-��&�da�t�-/��o�,�����i6��z�j�* A*\n���0e$��HH!B_Z3�k`�1�� m&2�7��2#������"�P���=!r�1t���Y�����ܪ+��V����T��ܖ5@z�Ӣ��+ʈ�;Yڎ}�Djעr����M^�H0A=R���P�Z�!�?�	jQ��ܡ���y���Ԛ���c�����&�`	y����ѹ�$3�Pm�r��
ђ��]�(6+�
������}'{�_W��n178���P��̀��ȉ��IqPpM���Fk-l|�[�g�Cń>f��+H��P��̢�U'>�-\�_�b����d��D)���C�-t4���֣��8@���+G���u���3��z8{����宑zꈞ����Q(�,��f�5H*�v(/2�R��X��MŞО�\�Z��<��7��7{�t.YnVQr/��4�Q�&+�'�����.�R��";xS���$��ܕ[�JI+���$���2eoY�#�((��}Z��X��\/ww�vPN��(2�?~������j���#u�&��b?��F�"�"��I�K��*��,Q��)�C�y��w���Y�0G����{*g�m���h�_����#F�Ȱ�r2���WX��wU?��^%k�J�q-��04{&��!" ?�Q QU�k"��B#dsȧ�u���zEHx���Ւ�1�M�H�ʂT�R�X�ki|�<���Y�5;��	��wuq���� 5��e.G�f���_-�S��!���k�����R%����0��P!���n��sP��%�C��=��5�a?����O���F��˦���%�߸`׿K�T��]�ŋ�,2������.pO�/��M/��A�hN�E"0�.�4Ձx�b�m�R`�eVT�`�K�JO>�R��P�0�I�^���@��t���xS���(��!���� îy����ާ��|���Q���@�'�{<��u[Q#�}eX��Օ��
���u�@�h�����S��>Կ&#l�תC�D�ڤ�gn��w�;�ǓH| k�����Z�O{��{�+�oǻ��ļ�>-��k�sZ]�u�ށO�̍�u���56t΍`,p�6ES�)�@�d�i�U�ʊ��?wO���n(�N	�ɏ�ώ�st$���v�ܝV�g���ɽ�����7?B	o�5��-�:=����I����=��y�2�8]D�NS�&� ��I
&>�iu�e
�.i��ƌPȳ�J�`��Ux1<fg�A��E��qFh`��x�!���6
�8���U��=�,o�	�b\�����M	"|H��O~��(��0�ͧXS��88���F�uUU J�@k�����K�P�x���ў)��.��:
���u�+�ˎ�E4�������Ƨ+u�U{4ц��%Qr�(�\ƽ�4�_�C��(��h7�@ƞ�3v�u�u SB����kT�:{m�5B�|<X�iWD+��sŠ�~n'�J�d4��p��5�~>�,P9o�8Ȃ�,�H�>��3Ὺx�J|Os�wY��vlsH#�d/�P����4~&�%	݌�(��d��D�I� �f�:�~X�Ra��3S����2y��zt˒|�yGS6e��J�+ń�<;����D?V�Nq�y��Q�P54����|�?�(�>��@��`�G6/x���t+ �9�9�uӁh}��?\HL��1?�߱�{"���	�ɉ�{=��m�H��r^��5����[;�>抰��!"S-�g%K�S�[�Ƨ�n�2�v)Li�* (�D"��������#���ɓd��	��iv�Ah�
�v�i�����</0W�܋�X*�8�멝�����䠋���J�?Ǔ����2�\�Ps7����R��*�/���4���_��s��&�I�R��s��(�r������H4��J6�S�iթ��Og78����z::N�0����2��}�>V3�R�̣��V���۹��uH�e�3�I>ʝm�H�MV3���OXp@�D�T�V��S�=��{��k������8pٟ\7��DY%,m�3+];�a[$F>WJ�O��)�D��S��e��0�YɷTu�vo��f��Ee
��&t��$�od�K�|�Po����1k���Vlt�}�3Q�
#�Dk�����^x���.֡�h�K�߇ڔmێ���:��)�\��p�g�l��n�܇Js����*����cw®̤�o���zc��K6��e�����h=��t3�UV�U�wK�c4H\��+9i�W%��Z�uy�9��$lҏ���ܼ��Vu�}2�*3��.���,�N�K;�Pr��B�l=����O��N�]��e���ѻ���s�ʿ����6��z�oȰy��_
:�3d�	�;Z�0�Q-��=G���^���;�X��A=������5Q�ƈ[�!�%���cy}�HeAC~�wºU���k��kآX3VL�p����W� �N�y��@�g4z�7x>���Bx�EG��oA��@gP�O�?=�<Ktd�Pũ��Q���K*
�Րs�M!X�e��0cc֪�Muùv���+e)�^ߏ�xuFԐ�V�������$F�uf6���%~�o��2����G�Fu�h��;.lz�����u�p3ab��cT���?*p�ɶ��$�|�$pwȕA��2�k�o��G�:�^ؼ�����`hmJ٭�ګ>����f���<b����c��&���k���C�	�7d��y�މI'*хV���VX�u���9k-JSJ=F��qI��y��uq���IOA/@I�3��U]�U/Y�2�GnR#`��߀�l���R��8E�ԟc�E1ݬ"�87�ò�o'�-Ґ�W��f9��_�fQ�W�t�V��y�q��7:w����K�I=Ɋ	89JN���g\��G֘3��ߧI�/�Q���8��	 �T�v9�8���?Nt��;�|7<�W�i��)5e�׎́+ ��2���eRmK��p,�7q��*��셅���u2����0Iȝ���I����G^uCs�<���S�:���f+D�I�o�~����=o�������`��>�aH?q��W�E�8]�o��o?�\a��R2��k���gt��Bf��}
�0+t�I�HO�r��(7h����u+c��ЈC�k\��ҋ���P���X��GSO tu|'�(���3�ld�A�zܝ�ln��(�4��:ܧ��Q<#>�gzՔ�I*Ʊ�Sn��G),y8�lA��Nq���ʡ_�L��bm�@DY�P}�l��$Z���^U=�_Y��i}`UK���?{�����ss�[1��`�Pt��쩜�Y;|����l^_N%^�P������٧V��Bb��e�{l`�mK1O��r�ӗ	n�)~��e��+��i�)×��q8#vMXq2�I���`��Υ�=�yihg�6�ށ9�#Q��XW�1�Lc��F�*I��vFDq<��Ŗ�4s��$�>S<�8������siF-CkEg$k��B'��,��K]2�෎�x�T�>����|r$�#�d��B�rV)���a>Mi#]��+�g�4i0a5��$ws{�����'����}�vApn��_:�b��!'�zz|�C�Bx��9=����f[y�t@c�J)pSnE���'�S�Z��5ɤ�@.buf�%�S���\�,μ�P��Z}3OY��=y��� 쌏�cl+�*�9�h��ܘ��dh	^|���b4]��1�S̫���ٻH��3�\��~�b��vo6�kL����OOwi���bQ�-G��s�?�qhuI4jv�xLs��������a��!��$��ř_�\;��,3�\�H�N�FܯmEC�ڃf��ڸ`ˉȏ�2I���#13��{�^0)�<�z@	���َ��gf��B�W�L���0�}�Ic�vn,�eA���{�d�"ϵ٫�H�ƺ�ԥ�j[� ��)6��b�"�R��p���ȡ���X��e��_wQ�k1%���Ŵ�y��mB��ۏ���۠f�w!� u �#Q��`�o�=s���ɺֺ�ݠ�d��8���A!�[�k���k/z�ܟ!�@���_��St���
5��7�`���bD+�Q8� 4v���E�-��h�=�ّڙ��E�UC4dd�f��F�hQ�����o�F-�1M�IV\�4ͱRu����
�Y�{3���O�,�m�[N��i�c$��N�THr�ǆc�zr�ۿ@��\1Nb_�0jhJ��ip���k�j�j*���έXi���pm�>�a��s����37���_w7������QƵ��Y�Y%����;��� cm�P@./�����>J/xj��$��^̰�+����
����B!�ub��`�-��9�t�кe��a�.��5�b{� v��Y��8eM��`l�<k����k%=�7>�\Z���3�^Ga��H�S���z�˞�_~����!�E{`��~8��̘�PF�� �s��Gf<U�@� *���M%�Ŀi�2�.�&��?;C�>�\��H���X��/ֳ�T�M�ed��`��z�L��9,�(�}�C�����~�6(_������=��{)t�P��gv���4k��g���"%e��`��Kts�ѫ��t�G�.񟗩Yf��y-)�����+�ot���ڍm�3)�*+���.�7v����\-N)�Yht�f��;U�"I��ڭB�!;��r�'��E�ʑ� QN����%�r!��2dTd�o��B��T����0e��7��(����)��&/B��]�����q�wB�B9?c�s϶�u��K5yn�:syi8S��(��D�������$+5]�X�@:�Ě��)��
8L��n��i1��X~
$C��{lC �|[�`�KH��W���n�#]:�,Nf��ZCS[��{��!IV�#��<��"�Bq�%,��h�^p샀��Q��h_o9C��l����� ��x_Q̹�
^a���ېU�.a�$҇�@W�I�2B��s>��Ӽ.�;|�c������Q!���K>2=��3�Wt��-Z�h��2�)w��	�ǣ}Dթ�5��G�	5̚�F��8�wA���`A��@~��*N��1�ΕC�O����F�>���x��:�-�7]>!���p�Ҽ�Wi����fSLut!FoojJl���BF�`�Vf������}�=!N������>�h΃����I����jw�f6T�uh�F��2�%(�
|�km�Zu��8���Mܯ��M�K�q	Q�Y�+���>rQ�)$�,�S+�1�EN�!ܙoy�Y�ڣ"5Ij|�*�=��Z�=�joG}2�?�4PB��Eg,K�:u��!Ν_��e�䢷���7��]K�<�i��	P���O;���]�册�D���ϑ*�=��9���J��+��V���d�
ڣ�}�8��4dV�r��Y��WA����	��-��}�|�>�[��T����7q6���f��o�(Y�绹v�S���-�����OFs`g���)�e9�S#&|� ~�n�u��1�#�����6��w�(�jG���Y,��I�V��nZصUı7�Q�&��\XV�Im><}!`Z�!�f �ǿ��x$/y��j�ŧ�~���]�\:�[��U�W�^&�N>pɝ�����7��YF|H�M�s��@F�ݳ��U���j��L��U0(��Y�1�6��{��N����Э�E��`�ړl�;{�㏜f�u��8����Va��
��I�,���F�>�t]=�c�N�u�AqM�)V�驔��	�K&��D��bWW"�����~F�[�Xn�.ƨ�o+�ݐ�h.H�:���$f�',��G�n�ƢCg�-N�[�|;�u�:�`36��h�j�n�GGB� M�'vx��]T��(eWJT��{�~L����:6���^n8`���yMc2���7-�H;��~ܭ+h.:�;>&���d�kǺ�_>�U~"�Q��O�*-�쮋�������Z��L�fZ�K�/l>�v�����ᨢ��ͭ�%$��M�H��О�2酛�C)��"��
M��<x�����M��ڏ��~5lS(�WT�}A��ę#�"�)�Y/@������%��t���� �3.&J�N����-�5��>�1�����=�6T�޸JU�^�4!��Y;7M#�6Gܸehǚ��A"}���qd���!V7^��X��h�MWIX�x�G_,.x{!55�9bW��Wb�Zϖ��'�2�=)Ή"����H���Э���R�P�R��:Q�����	�v�΂1�a�6�����F1��J��i�'�Y�$ߥX?3��{���-m��`�P]H���$ۘ�w`�Y�6�q.Ɯ?���q�2�#c
�����@n6�4���F���}A�CCs��hkix��z�%O�[�	��N����N�Z�-�����ncPAu�f��/��$�v���r�`���Lj26��[��Z-��}i����i5Qj+���%�����G)I�ӥ��bh��-V.yg!Kб�a�x�V|���'TX�l��-�+0)ʋ[Ρ�W��Z���)ZC�ǭ�"&��BCa�y\���-c#�~��&g(F.�[�g�29>�n��H#<���5��E���]�Ɍh� �N��v��~:�V�O�K�	�ϩ�3�����9��ҼgA�,����D\��Z���B�̴SrM��$4�I�a�� �����]e`��#�bw�L��+@�i_��$}�nj5e��p]��n���<o�b_^U,�%�EH�>��v���;w�uҀt2�ځ\�Z�Y�y�M�i��T�#�R@���� V?����0��~v��i�g=�����i��{]�d�</M�	�;�#J���U�V��Hq����G���"cqc=�+:pBɚ.}*�"'Y<d�X�� Ҧ�K"s��i�|����W���<�5�i�S�
�F�{f� ����y��jt O�b?�v�]�(�$h�rL��!�3Ӟ��4�%2�����T��k[B�2��QSF���K�#C�,���9"4=ʸ�h�)\��K�@�K|�4lީ�C5�1��:�i�h�{ 1ysN��E&��2Zڛ���㍧�#��09�U|��P)�3Xv����@��r4Iʳ�*z�ԣuv���c��u���.S�T�6�"+�n	k4��9�������_��%�$?x7���������}!#�J�LXK���8�u�?��t_��<�MROc��SҜ��~��Zx������6*��4�
���b�~��d�5���=�ڡ{��i��&��UJe�j-�w��[b��V��M��t ���� ~"�����cƳ�e}����yS��qyD_�䥌�I�Y�@�r�H�RO]T�<˂��FA��<)O��Y��e�wg s�^{���ܜ(���}\u�L`4ߤ�c��<�����Cv8���N��"��=#|#�g*mETB��_U�qg�=\��-���g������~�.Lc4}+�m�AR��f��mp��Hy�F��U��r��B8��[nCH���c��%ѧu�"<-�L�xe�=�o���l��UVBx���ҩ;��fռɆ�r��!p<���͗�/�b9�_���~��g�3o�89��	}��7̝]Ԙ���p
Of�����6{��/��Vq�?@F�l*Q�I��3��7 q�z���֡Z��ܠ�t����R�ԁXrH���_s�&���!���0��kݘ�Q%"g�?�+ɐ�o���d����u%��",����t�+�iq��H��p,�G����N��r�Z�d�h7_�wړN+��	ፒ^�W �x1��_f�lm�`5/d����e��rli��<�<���D^�F�uP#A)������+N*DB̓$�o�&;��YuW�oJ�����RpX�DD�=u�B6��V�Kb�_[2��A0�|��� 0���?�����s#DU�)M.�e��\�C�x�SgS��m��i���M�6��,<OP�ԡ'�ì�|6<0��B���4_�����ɟC��?��;�m�o����(6/��d�]���\hƝ������2nu@���	�W:�41�
 +��k��W{�-<�QVgy|Y��S��-m�c�
����c��dG���-awR��������ݒ8�����M�<��9��b;���!��T�`R�R�p-}2�t��2���$m�q>N2參��y��!m����%�;��`K�ʩd�T뇽�}�f��h�G�%��p��;�sY≪�	�ZzŦƚ(I�w{(ɖ������~����:�D���	;�@AA���-*�F��u��t�����.�����>������� �� �nh���?�P�!�&i��!J�|I���p4����w�2ܡ�2d�Uz��O/��W����"\H6�J0]��jQ�׮��s$Q��c��?v739r,�Yv��=�x<@ac+��~dh?��o4�~�N@-�-�M���$�$�jR��6�?�6z���@��������jh���
`�-�q��v�Q�5�0pC�d^�]�Nק!3t�9S\��%�>��.Ȋ���޼1Y���*�� ������V2�wk�WK�	�����E�t�E�>lT�����
`!P\�c������	m�8�ۯ� �5��
�Ak(SI3Ə���!�P���-��{�B��ϩ���o�%�9!�IF�\������Ò��z~o~4v{�B��s��E7#�A���Y������m�u�%�b��T�{�y�
[�󚱜�:f���$����1�܆�;�=T
X���>��a��������,P��В����$�r1&J�y�O�7j���3��,Qa?ᙥ�^�<:eoX�An�w;���s��L�}��&fKw�kCTπ���՗�ݏ�.�
�_��r�g���vo��1��'�W���ЫQF>	ǧ�C!Nf�)7ޗ; ,�n� WW��ǺbU���ܬ\�@}L��6���H!�Dw��A��p
�13ˮps�˰Q���b��#K:�H��Na�W�����z�p��A�m�R��'�O�\$U�Jm�^o9P�l��}A��yJ�y+\��j<>��;��\xW޺����?�	��j�;�H{��i�+�\,;Fg�4�rjTp_�蛸�&���SQHb�$���Q� œ\�W��o^~�!��F΄W�X�U5؈�!�ӷB�d�C,�� �T$}vf�pm@sv�2PN ��p�jeu��Hx�1��A�E��Ў���30̶�:���K��%����l[*���+2~�n��VG>N+_�`�C���u{����o��7~)���U��H���F����ĥ��c���]"�
�������~�-s]�}G$_�(\�8�&�Ij�G��vc�4�N��K�gs� Ji2��D�w�w�jR ��	9]�Yf��A��e=S��~Z�1�KaϘ5�k�o�u\Q�<v�qK����zE�����ǫB�1��p1S6QSM��h:�tXK^m޷j��?kϟ,�n���Z�I
4�MQ�bX�^;$H��f��o�;t�(,""iV���rFe|��jJ�9���\� �� /��L��R���	oah�k����G����=�}��P-�E �B�R7-E�����t5���x*�V�̻~Yh�B���_�R�R?�η&0BE?��ط��$o�茯9��n�g󙓘�K�$�4P&G�6���XQ��[��׌"�)a�M7�h W˺.>��-rT��߱u|@&j��l��S7s�������?Lޒ�����)�s�ٵv�)-�e]I�,�x9	������0�h"R��Jy[��m+~�n25��us̓��	trG2?�	�����o�~��9�?ٙKw� L��U
[�o�F k��Xqv���h��iGk�oB<_�;n���<!�/f�c��C���3�)?w�:#&�[`�䯆��|'�ڟ �q��L�΀}�ar��ѕ"o����c����f�D��-n�LriJ�[$S�X�!��_�$���ыNE���lA�2UúK�6�@���)����l��7oRi��(d���%�?>�dWutĨ?��؍H�<�fU��m��L�'����?�*귉-�����Q�G�J�)ֺno���)�fF��� ��M���֟��,l=���K��Enfs�i!�s�P��2���ǗU(����}������A]�0��^s|�s�%����s֡u\�_v�G�O�i�"J"�sl݉7�k~�Q-��èX��'�H^o�j��������i�\nK���DP�����W�
k�G1�L�5k3�b�c�t�/rn���g#1r���b����Ｓ�L *#?y>I
l�H� �ڊ\?��o`�E�\����&��Ɖ�g�!z��cn�ߑ.�%<�P/ܺ���-4�n	��,fÓ/��G�WF������}�^��y�3"�51��v'yp��>�힀-�TG�!26�C�"W5Sd��?���tyG۴rڪeC�5�ql)��}�S�u��]�ٻ�
h�z�V9Z���^�<e�V<�4��
y�l���<4�L�����(S�&E��h�#�XZ/�B�P��2"�h1'�]���h��").}9���)���P#е�H��2|,M�m�Sã�3l�>�Яʗ]���o���U��y� ��c�<���Ư�ur8����o~Cpus���^�4"{2b��x��+���D'QǏ���M���
$v���X�W%z�%;#�`�gp�\pU���$�l�$�`!�P�d�ղ�|�L�=�;�r٫\�<��ޤt�uq����2��������\�j3*]��f��0���������񢿧?�3~��Z��J�\t#�~�H��ߥ�A5���sV��#E�,�G�ũ{I��:ʰy���TQݶmn�� �����N�gҽ�<�7̕�n�lvk��iOv���圗���
mr���^�����,����"�*P%j�ñq��������)ȓ���@H�Ap{UHۂV��-٦�$�@D������kB��y�cǝ�7A�@�D�(��#�r�D%����<�C��3�ʾ~�qs=���n2��k�;D�q ��d��#Y�u�dD�-އ:��}bz�Y�׊i�	W]� +�G'?�����߰���h����_؃�l��j$�C��=wvB(�咏�x$=5���-�sV��PجԿ��wL_=8�?���ovkJ�6�=� )!�l?SS�������FAd�W��3&A��[������G�P	�dֹ��L�Cm��RպNTn}��a`$9h6�ڭ��&;(I����&�a	������WD?	�2�����6�O�Q�ȧ�����b6�\��Β���5�߱��X0\֤i*y�ʃ6C��R����
���m��6��W��ђ�d�@K	-��[�1����-��y�c �$��V��d��'R��9g��c��@<�+q3���s�4���{_�X�u�żW[6=K�&��`�K�\�N��֗��64�0*"Q=�>Z�{�0iA+�ui�k<�_�+㰦*&���f��b��hٚ)�%z��\�MP������Y���X�l���E���pc��i��4+�?}�*c�7�f�����]:)��{��vB枆]v�b�.��+��%�����禪'W�,D�� �xֱ��ȶ�D�${�="m��h<�K*3L�$J?z�_.fI��^�C���x�Q�}��� n�s�=�� �8���}nf���������ni�/�/O�L����DJ�n�E)��x�� Q�?���D�� �I�,�٠����������ߵg[Q�2�l�x�tR�sq芢�A��VD��G��Q����L�R��c)o�R�a{>��A�����A��f��h�]/K��`�BgT�~A���w�~M�K��n�/��$�TOd"�[s�܊|Dd8��2+=V���A8�*�%�e�hQ Ã���r!�|���\!�\R!t���V���P���6����	
OH%^aǈ5�!�ҹ{�c���#��<�6�O�;�"�����i�����i�LR�8�L�質M�A^��� Er��A*f(ޘ��;e��ݕ���س暡�Qq}����Ro��@��4R�-~��e���B�^_3p(��]�t�|S�M��o�6�w�i6v�I����NGtƫ{1l�O|^���u���J��'ί(%�NT�׈�8R���7w��V.{Qn�<�r�ȈsTlu�е����פֿ�����(�S9����o��
D��l��iE)t���� ?��^�� ��S1
�
+�L�^��FDh�6���x�S&�@pNZ�;�2�t�lǵU�V�~W�4� ���m��� jŉ����j;�g�
�_z�卺#T�:8���r^xK��<%�Tm>'����NV7�SZK���q��1>����o}�N\�Z��L�V�d��}kޟ��"�v=]_���,Cq�~�ˡ�i7�]�;�9�������F��R��)Io��YFK��A��3z���gj7�2�y�r*q��X�nu�Z�;OJ2!a�+,������Z����
RF�Y�~SG�dJJm��`m�:�ө��vP^�F(�w��g�r��P��k�YSIO�s#���G#�륪��WS��i2���O����W�i���^z�A �f㌝a���3��rsUՐY})�*/�X��[�2�M��O��,��'�w���16��d�G�@��6x&<$�1:���zt�~v:�L���R�+�		��Y�`�(Ya�X�!��dJZ,�tH?X���T7؉g�&�El�%)*8==��ר�k�V���z4�������c��N�*�t<≟��
#�>���`�ňn�T����S:�s\lO��m�����ӊ�J~A7n/�n�`iW�O,�=�jq����IW*���Y�_/���3+�(B_�)����2©V��C0�K[p)�bw��g��x����N|t?֍gD�������Of�<e���;kȍ�[���\�����D��wA�֟5�z+��6�$&��Ŭ�q<�)8��&"χ����	��K1Pݞ�䰨t\�M[�/��5g��}�P�n[���~����"+Ud�����D�u�2�5�#6gQ�<�
��� �7{���!����]�R(�J��X׮��JSխ�=���0�	�ȷ��E���h���B����Ns�aS�%�����a	����n��w�8~�$=�wY��F`�����t�@�p��cn�M�0fd�w�@�G�s�t �d����	q4���4&��gd�v�[G��n�0Z���x5ȝ�4�f!7�-�|UQ?
 $�+���� JF��	짼Ha��.Wg.̌�y�h��'f)d*@XU_�	V?��5f��y5\�D�A��4�dN��e���E���܆ŤA�ɋDl�hY�B���v=�<g���	djY^Uާ��W�E��g��mo���[5�p���H0��^��D7זZ������1ŀ��:ȃ�*���>�u��'��Z_@I��%(��n�\`���ɜ*T�ޤ�"�Q��1~mYy���beH���M�Q�o�w�Z>a;���F����cO���_� );��B04S��7|���zg��P��?�����U�~�ꦀ܎W>_��k%"��G���vg��DS3�35�u:�7K��x�ݕ)��2BՊ؏�fd��^@�OCL̬#���+�������_��SJ�;^+��c.d���k�	�JZW�a�NOE���� ^��'n2�F@*�z��.}ߥ \��4��%+U��g�P�h�K�-���[$ �����<�<r1���zV>�?��fֵhܾ@("P�8�"������*��p[j�#��W�'�h�˹А#L���	Mu�����iO*�ibMIe��Y��\�T�m�#�i�Ao)��n\�%�+~K�1w�`��&̞r	���S������(�
���l�<�Rz�j�#�<x�[��oLӯ�L��v�������6��7ӹ+��TnsL]���M�e�D���zL22�ܹ;�\y?�"��r��Q�w7�E�ONe�f�����9���Y��[9xR�Q&</F��I_���*�*�����󒋆�{�"��s��s�ޱ��q=�|��u�cH��=q�yJ����E~���S���W����w$>/���/ۜn�a�eb��J��a��|G���`ľ�M������;n%j8fz���#p�,�יU6��%�����w?+��m1�ɖ��������U#螋���ǭ�7R�8e���HXK(��_�P�N�=�E��� �1�"�:����v5c^�'^IJְ#��l3��U�λd�T*D1���E��D�;��3���3h/C&�o����M)aa~v���e!���^zR�V�����.:(*�[�m'/Z����u���A&�=3kKL�1z�S�>�ȭR����o��r�}���A��Z�^�I�x�/D	Y���������Ç���"��|��]�-u��i��F�t�.� �{�u����Z�b��4��b�'�\*
SV�de�Y B/��0�j�. ����O ���rQ{�'c�=�N���,â��}��Q� XCep�z��ڏE���B�V7ԩՑ�슕���G�C���+�w6��U���.�=k:���Z1%ޢ�L�uP�k@�����PcuZt~̢�������Qqhk-�����B�!�/�9L������dN�Dv6�����+oC��;m����:M��pn󚆜�0�u�Z��)�
�ʹ�cHݘ�lڼ��\A��9@���G1��h�r�՟�e���C �����Fv��CBN�G��3ZJBŁ#f��T��I��A?����)&Cqm�=���V�K.�7��5�v��uh�������w�iu��B�(�(�v����yS�"�j7���*2u�~�0�_x��~]��~E@�G�z�52M������ $�҂��;�F�>+���;��&t��X]ފq&�lv�n��œ���ƶ���o���*�F ީ{��J�S$�k���n�'�UQ�w������\(����j�_�F�}��^�?�X����;�w#�uo�`O2~9�L;��VJ~��3_&7�����9�O���-��U�u1�>=f̱� ��mr�d\0�4��=P>�;���3��{��`�����s�a5�ƲZ�R(�T�������1��l� l%�@:����E6���#eir��=��a0m��v����z�{3��nS���lչ�Z1� $�� �]g��vs�=�.$�ͽU8(1����c�U�����x���K�����'&���ֱ��|׌[�N�@M��a�/�%��NO������ʰ��s�e��
�~�Qv����5X��X}�pj#lFq"C��#p�5UR-�J#ni(�l��b��]4���'u�B���6ƤՀqБ��'�M�t��!��ߟ����#�3��+���q�"Z���ښ#A�����7$����O�q�0�r|����K�����o5��s�4L�n����Iop�+���;�a]��?Q<}pc�8��Z���/��b��3\���
�*���p�ɕY�Y/2x&���Ԋ��w�Qp����ێ���^5�X�Pa�4h�D������U(�԰��'�V���p���7�H���׬�M�-�����2.�^2��A�|1n7D��a����C��ߑ)�h�k�gM1@�˘W"�A��h��V�#JRm��
|��Gi/����3��IT�&q�������V��0�7����"���n[w�*�,� �y���#�;~Hed}���X:e�
��/��Y�}�f\��
Uޑ�J��7����1�Hм�?(�ڑ�v���V �_� z����}�ap���8e��&�aX�%� ��(K�Gn8bȜ�vu77��q/>�	�|��H��͘�WY��)Xi�"oFR�P��wgm
[� I�W�Sg���O�S>�S�d��v�"�01ڐ�v��� ����zo<e3?�{��E��Ђ̏�-C����"I���ZGA�(� mc�R�0�N�8���SkK�Og�z�ZS����[E��ʳت����{�N�--;P�*�L�pB�tB˽�~9�=M����OX�ab졚v?vyњ�FK�C�<K��~X�4��U@�O+���]�~���K���y%a�\�U2"'�7@��O� ���a�?bL(��1_�)g�8kt��g ǋ`�$c�e�W���r�ʻ�;ѥ2�3����j����}�U�lp�pP��Z	�f���[��_�@�=��O
�:�@�B�J�����*ߪi�	�+��N��o�%�g����Zx�vu�cS� >'iy�f.[��1��*�â5��(�bwV��8[
H�TW�P���tyJJ�_�I)�kb����P=�����L��WJ�䊡h�+��Հ�]�eݽ�(�@6v���k$�5�^z��U�(��2� r2E"y��md�7�|� Jmqe=1D�Ɇm�:�3�oq�8I��43�dj�v�LqX��-5E��Z���qP��D��R:�dK�����6!6�L�P���o��2�rH�"	\`�?>�i=vPS��mާ�M?��zjVj�6Z5N��n�C=�v��|��+�1���ط`�&��?fQK�zc�It�#�/t��H�V�[�Z��P�>�N�W����|��&��/��oԖ��䎶C��q<�f��2�d���y}-��Ȁ��R��5ig�wgK�4�m>_]�b�4�J��^����G��'����=օ���o�$I
�D��x<vٳ4 ��Ɩn�LR��X�kl��ʲ9��<�*@��PԼc��@�����%�\�f��pĨ�;Zw�`B�Q�P>�<�l�J8�0�B�顮N:���3r�0^-��@�=G��dy�Vo����@l��E"�fj@��]?��Y		��-�&�I�hl%�����+ԃ�̖�«�q�]'��mW�)a�bN��f��P�$�*P]J��ψ�$3������09q���=宴PV�]ڂ��NnKC9f%�g��=���A������w�EY�pJ�;�1��+$�,�~le���<��G���.�6vDM������=n���LP��	{d����uT:q�]D�E�����=l1"��������v^���4n��Q��2��#- \~��|K{�Z�/�#M�O�c�| ��_�����vd�-���8yEk��#�-+V�2/�N��|ͼ��JS��D�:BG镔�11�YJ���4˞ぬ,�L�>�`�w�8UUl�Uu��On����W����֭9B�%.;Ć��Q��CI�v<l�{O&�@@��r�.u�a@;�S��]��.��7zգ���ΘFw����g�h��n,���1�:���P�s!c�����Ԥ�]���V�='޻�'�I�vw��Rȗn�Og[Ҿm�^	�����+��r�s��X)٪�T��"1��iʆa�+���~�iz8Uнmf�"�+��9�<0�8�
���g	d�����v#c6l��+����M��絤�ü�I�!)[������'����qH��`�Z����`i;��+�N��}OsS��O�RnP��r��zN4jh��d���(0��JW�I�v�����G�w$G\�Q���8�G��EfP�Dx=+ٽ4�-��f��M�-/t&��mX>w�������_(��%�Ip��j���e���JY��)]�v^�/���ZAO�o+*rؾ_ >g��kNBkX5f�帢��UW���J����eS���{�r!��$�����loLt���0ol��J\ p�u)JZj}�!ȍh�(X�B(�S��Meh��E��i�fV=�Z6HĊ��3��c0�����ͿE<�VA�ﺧ�kݔ+�{�*��8�b�=�J �y��Ǜ�6$"�["�W;Cz�qa�oM���djϾ�����]����y8�ys����Za��gM�Y�
S<{�22�5��E�
}� �3�HF��uNV;q��3EH��$h�����G���Sօ�(j��K�Ry\0��N�.Q��c�`C�r\��q���-1��k���H�.ص����w�*��O��������ʼ�23Y�����܊���R�Ѽ�&Q��G���QX\��LXe$ӊ��	-� ��үEÂ8$dQy����|�n�|z�*_��"�3ZGC�F�Ϟ+*;+�I�!�om��b����z:�PW
A� �X�+@�?��yM��dS�Y�q-��hR�f�7m��\twz��-�Z��Rp���!O묟*�߶�m
u������9\�Q
Ax^�T���e�A�mfR���΍u�Ҡobh���L����֋�KhNE���=G$�m{��vG������Y�u���m��fȼ�N;gC����䷛�.����s�/�B�@�� :{N^�m��Ņ��\�g!����ZI�[%��"���x����C1z��~��=X�V0�2���7D��O{�9s!o ���5�3����l.ڀ�0�W��1�L:K�c&����&��é��?l���tIY�|����1� �^(F�Ѧ������:T]��R���Ԟ%��J��[2Z�Uuz�%�l� @d��F��9���P�a/v��!�1\���؃�5M��mq�ڿ�nਉ~Z�����o�����������	�$�^8��/�<�$���N��u�(���v��Lr��E7�~b�_/h���g���H��#��E|�x���ΊcY}P�ާ;�x�d�z	�:�&��N0U��0������#K�5��d��֝*j��H��Q�P�+"�����k�th�3z�kF��{���VB�L�TL����@�H�0@��	O`��� nh#[��O2ލ���.���(9���!r�r�� S��`D�&?A4$j�'+�L��ltQ(CwD�,>�#kg�l�5��a��9����o�Y�A���`�X���qZ�͕E���!��xT���5K�t�[��r�@�<��`�_�u�2iڝ���R�p0���Y̾��$���9�^��B> �;l�lL/��I�5o��AS�ҷ��-	���Pz�&(��I2wi/��?��/�R�n�~�ZF�}c�2�^��t#�*2��48P�!��F�`��g��&���|��_̘��l�ȸfYG�E�g@C�y�Q� �Cb�>���$�u2�nNBMf �93\Z�<R�~L�Z��A���)~E����S��Ӄu��M��J����xr����׶�g�DP�W$LݥK�M��	�\w��M?�rt��)�:e�Z�	�$l��.���U���)�����G�������4�B�aQ7�Rs�܅�
�t������G�� ;�1���V*��NZ/�}c3��ni�:O�Q}R��|�j�v�c��������5SC��t�=�|ޯ�'�K�)߶��G��}��_����ޅ�Z����Qg�9����v��<��j�,-�Y�\QO���@:��b!�D��-Q��(Pt��4�Ctw6��V��nӧ#���c��ccG�<<URH$x�r��E#"3������Dʉ�����ʨ[��ØB��kX(��K
�l���{�y������s�}̃3�a/��_2t*���c�5|��׸�Ђ�i�����?��Iҵ��A�&Fĥ�����33]���©�f3�1���μ>Y���C�ڋ�q:B��;�F��S��пg-�լT��~e�b
�4��<��G<-K�E�:z�w}-?�
<�ޜ���g�gi���pǪ���}�W#W�	�}��:�k��&���x�VG¶<K���Dkx��?i�S�� ����x8-ż$}��u�dY�	D�<] ��<�����J�4�a~L�O��&�k�3�jͿ��V9N�c����ţ-6��G���^� *�&�>T�g�ĲQ�&���]���Lhbf?	¨���[��?�)"��E'5L�� y��c��?��� ��,���H��#����fW�_��POU���c��d���)��`Ǘ�q�M���`��:��N�Үk���K�����z����@e�x���A��`�4��.c�Dkz�=�H�l��>3!U�W+�]�v��L����MB<V��#��=�@�"�t.mA��<����G���C��V�YY~�I:ԧ2;~g|E��T�[P�������f��>��*�W�+�;#	��^��pB���c}r��ɇ�"�'�{م�\�Pg�����FBZ��W�L���)���1Gt�)�^;�|�y���Y�Q�Jm`A��ÎM��a&x���Üu�gȘ�9��;��N��u�,FVe�q����]�-�1��|@�)6X(A���}�Ԁ
�pi���ߝ,�J�<D�3y�\"d�i]�U&���2
;j��žPП4�_�[�Vĵ%���#��Kp,c��3��#st0�g�Aa�N�t�y���K	���@��4K���M��s>34�x}*�"k�-��Q`���z�bjMo.�`J�PY�|����Sߛ�3�|wD�dR O�<_��)]���̔����aC֫N/g��-�\�~4ā��hS�k��a�t�YdJ�~ս7�$����Ά�'�5U	�.��\����H<R+������d�s�'<ot�'�3�gH:0��'�fU|��K6ym��l�w
Ȑ�=T��蝽����2S1"F	 U�Wy?JwI���N;���Q��/�*�a�l�W^�	b��3�{챰� ^�;S�#��" ȯ{���������~k�2���yx1��Hh�V%�R��+@E)�x�F)����ݮ$iX}Η������z�0�k��ߊu)ns|.��
���A#�;l�ׯ��|D��L;o����|W_���:S�=����0������ݤ>���;�A93�!��E�����)�+)�B�� ����tY\ ��K�0�݉x�{[��R����GH�e��▰i(|�H�_3��Q�;�ht)THq�`>$1x��B�%ֵ/��F�4�h��g�V��Ñ<�[�j�5�`�<���bR�4���P���&~1�������|�֊�y�J��m�^���'eޕ� +ڧ�\�n4�R�pzɍ��+4KAbWS��}��Ջ�R�k�\���L���,��H ����>"��J��}���k�f�BVv�+C���z<�y�R7��g���:��'7���#9Lf�a��Ġ$��Ư��+�^�p� <n��6�DE�-��k���<c��K1�>��7D�襅*&�W�Z�hD��x7����	:4|�Y�4��S��@8@z"�ׅ�N+f@p\���t�č�����i��S��l#� �i�x�;�������U9���ߵ�Xs��+v�V��w���g����JǴ�L��jw`�ȝ��;�7{��g7��k��^�H�4���)���.�b�亪hnc����
b+j&�ˬ̂�wu��:d���
@�����(
��ƑǤ��b����r�Sm�BZ�8.�fGί�jA?�;qW]�,�u,mϾc�z?I���kO�	U����p R|(���-���q�{5�:�FOFa٥o�~��DScFZba���,n�9ۤm�鷳�|g������U�%H}Z4�ޕ�yL���d۸�>���T A���4W-l��|�@���z.Eyᡶio��O)�#�_l��}��Í�FώY��tMr&��2�����Q%��ą�h���²��������e�s��-`����1���t����4��Վ]%�����1�����J��~Y�[��?t�Ҵ�^����4)�O�ϸ�R6����U�`��Ƃ�d���$R��Du�b|%��`���+�	R�zx��Z.��!d�C�SY�qR��A��X�`���6���^	�;U OE$.�1 bW]/
]s����OFV@���,����zKwZk-b���s����D�9_�]�$?�m�j�ӆ=K@��D1�c���aĵ��_��K"P�%GV�h6H8��ҵ���瀯�۳�4Ӣ~;1�|۩�;@��n�f|��tvT�A3��Y7�cn�=�nw�>����2;m�w5�&�
��@]E#�}~��+8D�N�5ܶm���̌�<X�R�jTA�d�����*��ՀF�;F�����kH)o����e� k蹴1OB/�^o;��k�����ę,
����N"
<�RknNi�#���L�Sb�ng���(.����\X:6�Tt���J}ew�m���-*�(������Dݮ�(� �>�bೊ#�6jH�"�Ybao�� �k&N�5^Է��ŵ��YZ��`T�^�q��ƟB��d=�T�:�d����H.�?cN�/�nDH�a4F���cr1O)�{��O�п�����d�ȅ�V����R�+϶��<�D���U��T<C�� ��71��O��XPc�n�Ey6t�	gߗ̷���ƨ8?�1+͌�
�� 6ܙ�s}t����}����s�{0��N�i�u4]n3��Ƀ�}x
��y�O�g��
�@3n�g�FEDR�'�_�8M�v��?2[������~��}��!���?"��w����A �����W\�K!f��oHs7���4��� �-��5���	fa�ᾝm�D�g"z\�߬��:/�f�����׆�y�����8���X����L�.Ъ�h�	��>�U`v��@�FZ\���i7��,��(��5tN^n�̙.+��o������� c��E3]p����`�6�J��(��8��+!Wsz��gK�B�����zX�A qZ�-�Ǔ�H!f�b���6�'z�������,c(�P'�8 )W�7;e��gGV8��>h�0[S�Ǫb4w�Q0��)cW.rq�޷�B�DŰ4K�̦{��O\`�'D��q�`k���?�g���/g�׋��>��p��T�2+Xs�9�����S��z��mJ7u��>��ᣪ�z���FW(�Hdc�'�V\��j�2�X#Ɔx�.�-o�O��DX[� i��m��	�O��%�Ǝѯ�.��U�uyPaėLCZS�_}%�j���mj.�L ��y��>d�\���T�n���r7V��7��G�kmD"׳��3y>��ы/�;��&�����IO�+?z���iG*��y�Ibu���+����S��P:�6Y�dx�2�����W�?� ��&�ţ��B�յ���X*勺<�Xv-�����G�+oKφ�C�0@i�_�u�����s��s�5�������L�lʂ;X@:b2'9k�Q�᾽�)"D�H��ܶ��Y�u;�����f�\T��ߴbV|na8���ޙmE�Y�(c�Ӑ�m+{֥�m�k�8���)6��;@(3~�'�q�X��7O��4@*��ӕn��5��Uȗ	!r��֐&�%^�A	�:{<�cGŶ��F�`FHY��U��s t���*Ɖ�i���3��^D=@-���@��Caz��?��l6�^d����ok�s���T�}g������}�i��m�M�o�`�"2���}���N�٬�����:Y�K���m�(����܄_k9ݰD2����=��*h���m��!E��p��>�j��z}Ke�b�}/�Y�m��g���├�9�,\*�Q�N�̕GQHr[=��_(�T��T�9�$�1~a0�Fa"#dY�\�cw��X�L�=u��}� �E�^�q���E�<ݢ�|������X�ָ/h��@��)rR���*��]���^���l D�<�RL�N�9�>����'�hK
kw����A*�C&���!y ��c��m��$>��I$T{�6�R�<�P�\]��͘���49�v`5sB(��g�￝l̀i�K���e�=��ge���Q�5��j9.�~(8���W$O���=��˧��x�Z�]4���[���R��L����U²O�:T��+c�|uy ��ڱ1������'�]���<J�p�0|��H�k��.�]��ZP�aʼ��Ys�bH�ZzO���~ ��ط2��4Z�4\�U$L�}%��Ĝ��({Zq�L��p,��ܤ���@���%���@^H���$&	JSr�n��������V,)����Ͽ��Η�[����z4�&��GFQB��X4�j}hQ��-�uے	MuQ�H*���O�m�l}�B����O�ŋ=�=�Ky���ϥ��j��|*���ײ�tǞ���}/i�,�'��I�U�T��/�O�S餴~<&@[���a0�=������k�f�~Z����8΋Rb*�}�r ���*�ڰ��'%����mu��<LG���G��І֙h�Qfފ�ܠ�[�
-)L�;��TV	Z��[ֲd.=g�{]���PQ��&Yw'u�-m�*qA>�T��#�Y�:�.n�~.��#I��*�:C�]�@jb?4�b��;12Vj2Ct��� .Y������!_�d���E���&�Yt�Ζ�.X�zD���������%�d��s��6�����'�5āT�w�]ڵ�����<�|S+�۴�B)dΥ+���'KgJ���@K��#�T|0��[AF�Q9��:�1��
7 (k�T��a�{�$嬆��&d�S(��p�~To�!�k�ޜx���@c�.�qg�ah$0��`4�����x�VQ�j��E:�Oؔ�Y-9G�8��K�!��Z�!����Kw�*"~�Ŭ��AR��
�	j*�3��b^�͡>����~o���e��Q>b��j�k3&������q���>�H�*��-�p+Y�j[�A�SI�I�յs���R�5�I��BĦv"��mLʁ��>�*>���_�����;su�����i�|�'r���������(��KP7%^�
F�Ľ:lDMDg�������I[�*:��t{C3�5���W�l����̦��G�#��`�B���r�N;�Yyv�>���/-IYg�<��ò����Yn���L"����Wyw �KM��P��c	gR&�zY,m`��/�&?�����@;��� ��`U�9�I&�ִ3��ђ�^@.8/�i�mt�!Z/����=9������+�`P&hәk�Oj���8�L�����n�����zi��D $�-�ʻh�{	�[Y�W�hz�y���мHP�a���-�A�1-��oz!���k]��mChD}6+-����)SU޶����!F�u��8�K�!�:�>RVh�����J�/����"d$�r?}ꥅ���J�g���/��;�F�͖�B>����4�� YU6�i�b§%}o�a�7=������W�իK��
}  }�����t��V56q>�~��a���p�,����g�L���E��ɋ�'���t����r�v[Ā�VR*�+�'�$�s�t�ӯ��\���Y���u��h�dnbu-��V�nw��D���N��0~҂�m+�t3-0]x�_ͅ�ܞF�s��l���y
�r�a�¥.���!E�Q�j��c��  ܿ�|g�0f�G/&��Vǉ��Ov8Lo)8�9jl�"���
���]M��Ɇ7wa�'��~s~X���L��؂��Q�O������MN
|%��� p ���P����ف�b��+D�yH��[)4t��x9;(�����I�"b����QV�_~�k'��bV�E4t�J��-��92��V�������$���"���sJ�E�|���71��Pb:X�����V����-�D�dҙ�s�l�������@U��ezG�k� `��V���]�L3�ܛ�V���WZ$ir���:~��*3���k�9�&�$麐X~�'��y�H�R�Tω�TK'���:-sH�P$�3��Ȕ/j�N�״��A��FMW�߷!2O�YB��q����c�P���2���}��.��R&��lpG�@�X�i1N�9�T����:�xH9!�:�Lk�����L�+f�r
����*=������t(� ~�"��>d���ܴ&�����mg�
Ô��x�&��kb�C��׶�j���N��
�D$����;#C%Da.�@v�n�Ñ���X�2zsq��|�?{.,��t��c0��
X�l���9rd�� �(��KмԺ����[�'o�d=e���/ ڟ�WT>59�j���+ �y"	5D[�w���}�E"&�S�M5u�cf{$J�Wb/|��p���d*���}��"�x�9fh,�y���!klw���
?��b�3��F6 @�1֜�_	
x�&`5�ՉPXz��=�~�ە���f�%�xS�3��+%�,���h�+�D=�D�v
YβTE��[Ym&�aj��.AӸ��]�b����!��U ��	��#L��|�ӵC:����MP �<J�3P�aF-ٮ��[ٕ�7�= �4���hCO�>v��2�7^�@�����g@�W���㹧(Ae���O�$��S.9?��D�Ϲ1����v?W ]59���&�W#��%Pb��L Љ��ž2���7k��z�<s*�>��ӈl+�cIo�sLKyX\i9�t(igCH�G��ѻ8�~>�O�
��Ek�֦�,k���5�t�x�)۳�� Mmb�)�Ծ�OXґ��#]8��w�kW��s�B�T�u���?1�oH� ڸ[~���T�OZ��ar���Ċh��O�8��+���i�j�%*��צ�q���0��ڔO�&��q�6���lsl_�$�s���=$�)e�|qr�[�/�W/�D�niM}Z�����n&��'�ÚH�l~�#���i�0+��H�w�܅�̜I���͆(ē2�N���\̀<��pGx��g����������T=i�eY���~ٗ��YM3�r������P"��8�����л����B�"�i`��d��+���f�}9폻��u�WȞ���#n�4Ɩ^�b�(���S<o�1н"����:�2�ħ�?��������4�Sg>C�]���Lr��U~Юy���`c9��Xo �W�/�L�ʸ������t���W���m�9u���6�E�Fw̖���۟��N�z=HR0B��>!L��U�&*2&��"L��Q���[�>M=k���o 災2b�ג�-�=2v�յŽE�-W[b��=�2����@#$�����Y�y�L+�$�8��G�;q�(I�`�R,:��-��G	ۣ�NIƾ��-J��l�Ԅ��٧U�=�i.�D9�+̀(��jUM��W�h>�x��l⋽L�a�2���nWB]ZT�9��OՈKS��K���]�"���O��L�ٟ1�Gizk��ֹ����s�(��j�`3y���Qo�������H�Q����u7�,���w�9�L*>���9M����Z­��A�DC��ޙ|��*J"������d�t 찣��i��rG�����i�n�u�0x��o1���P'�ݿ�9"��&2;��_u9Cs)���A*�`x�������^u����?��Ǡ��rƋ'���6��Bf�gCr+�!5!�N�fN�K��I�"��}U
ky�6x�fAҨ\��X���.��̃b�%+��u�n�h�w�l?G*����')
��Js`��}� \b&Ei��SZ�wc��8�5��t�RUzOn�4mx
�3+�������p���p�YS�c��2���|��}gCb΀�*q@e�m�&O8�ag̙,Ym��̶|��̴%������~ΐ�A]��r�Aʤ������v,�XI���[����Dj��]Z8���(��y�r����M̦��6.�nׯin�w[��Dk�2a��^�/��t����]���I��[ϋ>��c2���Q��h�ܠ��2���o��d��1|:ҫM��L�SܼC���:��TX��5�2$�N:�h�؎Q��M���Wjp�8��EI�'/q=�Y��2������'H�YOX�a��nC[8�ԣ ��֬h>�,�o�����س��?8���,\,�_������έ�mc�y^;��wh��*����G���9�y�uň��[��M#�qֈ���黽}>*�&W��i��	���_�U7؝��5>��c���t��+��NPc
o�7Pɐ�ρ/���� �-�:�]�Xd[V�w3W@Þ� ������^ ���ۺE�����\�P��z�`�st���#I�t�;�M�X�1>5�L���9�����OZ�~�H;q[�ߥ�
�\�Bh�v��fE��F:���~��v V?��6n%�$�0gF[���O����C���c�/J��S�s�X;�G�ؾx�M�?��IL���F)�	ȑR��~ 5}�D��a�������33?t+��CL�ypj�Nᯌ��r������W$�Fwy=	� 5�K���'l�;ۄ��P_C����yi	}I�H��9��[��@��Ώ�1ڀp),R�����j�
٣�W�^��l&2��s4�������Q�����0�]��Vz�H�}��	Z�ds݊�z.P�#�J�[|��n���L�O�6���7�}�|��z� �;��"�pb)
6� $�/����m�-�l�;w�(-��\#-�:Є���g2�3<�@`q�g� ֔%�36�f��}h m�1<~̥�+�Rn?7x%�u��-X��]�d�� ���n-�M������r0�����j����!bm��6A�v�Fߟ˂���Ӡ�3e���w����:{``�d���ȃU�[�#�� ::�|Fj r'�=�,�(D C�pk�
C��<�-�E�uՖ|M4O��B6	����y��F���,Q��8M<_�ype>��9�=����@D�����@��a�!���ӕ�a׆�ȟk/��[�a���S�I	�H����o7�����wQ˫<P��<�����a6�p�r�wF�9�	�~�_��U��" ��6?�8uOI�Z@�T��3���[��f+8@�l�3�5�o�������$�`�̗����y��I)��B!l���fy>h@��`��u[S��1���l���5G5���4K~��"Ć�L�G�c��rT���W)#�N�����'x����"�h����<��;9i�ذ��<��V��6��Cj{���&4t���X�1_2$�-H�Ģe}xe2�|��f�*��s�� �Њ�!��O�
��?�	ϭ"M�OF`�q�B��7׼H���W�o��XGF5����!�Rz%Wt����S��I��7_�����)���"/����5���tJ"�FJw�(ńIY�WG'�0^E���"wthgZ(H�?���3��"^��GD�?6i5BEn_��Xlq��a�K���Ek|����Soc�+�>�5��&������\�)I߾�pH40�r�,m�ϊ\,���DiB ���0&OaA��ٓ!���$��{x�&O���0���iO��n��oO�uir��quY��˂�^�yO�Պ�/xec���W��!�}z&��k��nY������`=�r7�^�i�|vW$C&�H�,Hn<��#IMU��EQ`h{ ����;�r5���!b�\�Bqʼ������,��_I$Kr꣱��-�Wsx%De��)/�t���ь6�� &5�sq��`[�CAPqv�����Ï�9A\bG59�꞊1�����֬���j�}nZYt	B�M��e�"�x��/�K�ӑ_&}�ի��阕2��<�OS)账�}M>C���1�N��+(7с�N�b�B�8�ϑVX����]X�v;v��F���9��q�_��\"�7 ^J�U[6h�=�V��|ގ�08�/��WE0sGF�oL�%�+�q/$�;��[���H��s�Zg1|y]"�?��d�$:xސ|��O�N0<���/pxUޣ���=UC��']�@�00��wѷ�!�h��62[�$fGcj�
���m>����X�����!�������"�Tm��Z����}.�J���2?��-�[Ӌ4�,x�j2y����$��n�MӤ��2�D�;�i�1,a�>��ǘ�-�I�y�*e��,� m��.Q;���^��9����%���ׂG��x�s� ������!�����q�.��B��p9�B��4�j��1A���� �ϱ��j��.��|��i�"4�.c���}��M?��������+yU��r����Ҡ�3�nh?=9�l=6Q�0+�����\\	!(MT#���$LZ���A*VC�b��~�\sr���ȕ����*
o��vL��`��!���Ѩ�pgCX�>'�_���D>�!�Y��;q���j���J\���pg���w6����|`����?�?�Z�;ȏ������Ȯ��|fd�J=���{��)���}��3{�]��\���dP�sϿ� ��2#�Zº�L�an��^��`�9�����Ƹ�:����O��<a&��\�����r��Z�� 0�@�@"�^���8�
1Cb?ZuP��Z�~�$�o�)A]�#YV�U5K���v�2�-}����,v!:	3�!aíD:v`n�d�pRT��&ڒ6���*P`�"{П��hy�qGb Z2�n�14��4��}j=��k��W���?�]�[75���\��o�Z�a���}�B�^�e�����.K�궂���.��C�?��u���H�㽯E>��d�_�_��R%ʍ�JQ�Dj߱�n��̱�������D]���<Ч,�Aw�s�Z�����}�>�S��rl5��9�+����\��'z���	v'ԥ�-�oÑ�`�����XT���v��Vg����rR}W\�=L������c���"h}�@����&7�n_D�ј~+A��Ṙ�y�����	�8&EL��'J뾿xh�I�.�b�r���v�>7�a��1V�4A^K1���x3�6�H+�l�m��3�0㏯���y@x��*�=�:��-=A}K]A��X��5�J����=�e���q�Yl)$��c
R&Yl�����괁O@��h�BH<CY�>.*^�f5B�j�/)�!��G�3ʋ��{�^��C�8��@�\�&lȖt ���/
� rw%-]����u	�q�6O-nT%��7�8{���TƱ�@D`�������?[�J���O�A�Rk.�ͯ�p�]P��q��B����k��y��tv%��=���uc�!��-:��D��s��L�����~|��AqS��`
~p�
r�/����4��ogRXaaMDw�b�T~wq0G>~����.\/����>�j��b�_Pc��BL�@�������.ɠ��jjp(7g��C-���M�6M�MѩIF�~�	'4َ0R�PĆ?+c�?�@���Ab�!��i�i����I���k��826YŶ�:r�
���/Kc�2`!��ٚ7�ˀc�3������8�_q=�ΐ��PD,��h?S^�O�x�]�糨�t�q��q�����1f��M,m��A�x��b�Y��*WFmGt�@e6ތ�i�ct����X��z��C�����H�ɛ�\���b�\�(�(Q�xG�3t?.з0�Bl�y0ψ#ẹ˪�Lv_hh��u���'[�-������r$�,������A��u�`M��a\������L����ʏ84�pKcgN�'OM��XEv�+��,43��������С]�:\����Oh���Y�2k�<�0��#��.%,\��1�"WK�p���7���h*�J(.��Ү�g�(�P 㟳�S�X�`�0-PB��S��\d���P��z�X�I��>��f��+NX�#"˞?I2�P�MA>�	�'6۵/J�\�T^ ����zD��oHS�^��tO-�teɎ|C�������Tϰ�!��b8���7y�ǜ$a�{�P�eC�7h�V4����o4%fZ�Z��h��"�Y�A����q�RI��Kts\<���Ŝ@L55-l��Bj���,C�Ģ�U�3H��v���`|:�\�S*?�t����G|�ŉ��I�f��%�7���Yf5��rv�C��s�1A����$v)c�Ob� �F��]:=���(�7 �h��@�.D�ʽ�Tի>�ז�J�)���#W�}�p�ce��a7U�2v�E�B�SZ开a�ޮ*����eg|>a����#X�6Ю�K�,�P��D�W����Tt� hZ��7Zq[���;O���|�C�� �fb)�p��-�e^��S.��Da���LO�v��j��C��x1{7i\�TE�$���B &����lBG�2��������XBIPs�%h�6�����"���]��VȽ]G�b��}J[Z}̓L�o�`��_���CY�0�P�Cr�%_Z����k������@�,��D���<r��k�H�x�梶zqqJ�������!��r.�#�9y��s�4U]�o�y��������4=��^cwuf�����D@�LclD��z5M��A~�c��K�a����a�X�4CT2�jz�HƠ�ͭ��|��|�)/y61JK
B�uP�$7%��<U�]⠆]�HI�3/�ig��`O��%6���Hl�����.��r!�ꝵ+'/���.��7�}��k}�I�T&���@d�~�l�EjFj� ?SISb�������?EѼ�N�����[�\=k�X�pIG=;�ڡ���u-S�#�e�?�����6؜��Ҁ�ƿ����cY��� ��Z[Y[��s2zzq�ރ��\k�_J�ٱ���.�"���~��ܜ�@T1����;N�x{|�p�p׭��Q�5��h����������fJ��m�~�,��#U�k�ZC�E�#R'�?,'F���y�.�|�ӻ�|�J�� B�� KQJl(��-��#Q�qq�E���ZUz�ß�=7_�L��=�\S�M3�I{�1�H�����b-�6�9���ց�j�\�����۟�d����q~�Ā�'�/T�8mY[�8�
>���;�<}�@ 1�q�rH���-GT��(��dM�u���Hr�������(c�"1Ktͧ�*�%���T%�cr`��������ݦ�wh9�|g�Z�`�3"�?X���V٨�B������q:�KqؔOeB�XL�]w��ٟME۟�Br��b���4,��uU��5*IB
UJ:�����8D*��;��w�l=����Ҳ�� ��b���a>sj�_�|V�#^ ���/��C<�����߃�(҂qp�C�=]�6;��=��ؔ�7a���j���ZQА�J	��N�_��%�ᘆ�,��u�9��g%Z��W\�D{~v�T���3�j	��dQ�5Y׸a�:�,���#t��(Lj��Y�ϼ���q�� �/ղk�lsɇ���AwJw&�_���7�ݙ�n6��>CN�F���B�I�{V�����:)  -��d�A��)�I�0y0��׃'6�����ϴ���YI��Ӗ�[V�_a�6U�YZ��Ț"�'ڐ���g�n�Ed�X�֫z[JU��s�%���%q�n��`�=#K���hG�v�"
��IE�e������`��A��[���!�����?\GL�.���_
�fI��=�*B��I������ݜ>�}»��|
�rZ�g����f_���Y�Zp����vֆ@�;�y����wx6?9>�na��hi�b�P2���|�R҈���E�+�P�W����=Ny�)��6��'E3ف��qm&R�%dqȾ'ԩ��ubx*���O?�^�.H�1Ô�#(�����[c��N�������W�o���'UG�����Z�<L�{�*ލ6�J���\��]CȤ�I�|~�D���=�����ʩ�ŗV%�J�!ȫ���)���L��J,.]`�$���I���
U�)܇����5�{Dk6&��Q��[i8k�9זy�q�L!Ĺ(�N���ڻ���);�*^���J5uţ���,��;K�E�	W���e�}���~/T�yE��k�o��,[;*�����	�� y���},��xD��T��O�8N�!M{yI�M�Q�{a��Y�A@�Խ�&1�du���Z�Boy�` �D�E��(�G&�ć�.�p���0O�)W���'D$�2~���t�|�*H���:s�`�v�c4"��  ���>��{��!8�HΨ߲�\8əc�z�o��c�������e܌��Al��B�0Nl�Dq>GL����YQ��Ǧhv�}�_�ɵ�sڟ9���]E��,�[M�ʶ%�cQyw��a�H�����B��@`�2'9����Q���Y�JK3��&����KL�[��G�����>[ŵ� w��n�t�ྫྷ��hv{�X�V[�o�jw$�i��ډ֑�.��+VgGq��yP*	�o���Q1q�L�Lw�/R�`��Y��\���V(���=�2�9���3�{������B�;!�%���D7o���E���bX�
�4�y���?C��Y��N�"��a`jW�1�a �EVH��v�_��nVk`0��:{���K�Zɼ�i?�
k���f��Ai�庨�Q�D�y��������*]�h�m�\ ���[�d^���p�7<�}�,HH�`ʶt�n�Yg#&���7���^��5��b���9g�}����*.
O[5��ItVKE��X�G�`-\h���gBݸŁ�/����b�,)��j��iq��P̬�s|Z�ka�WSǜ~��꟨��M汝��R	�l�IݗQ~< ��_ꔖ�̚�!fXE��\�����FbID��h{��C=3{���.�k��Ժy
H�/�]�mY��P��zRjOG�Aoo�4e�L^��x{!K �h��lk6"f�lQck���<
$q}X��d�����-��4��M%ڎi�t�R�P�����+d�o�Q9�� "��������{v�XJ1���4����g#y͌kO��VLd��B����������U�;�sz��o������+w��}D��X�5�2��Ҫ�&W�')ᙻ%����C�'rS���ا��������#P�{�$����d���V]�F�-u��*�N6�.�z&H�H��xʽR+�2G�T:�k<L��̏���|��{J��.��a-�?S��۷�3�hT��_f��U�$	�~+����$��4U5���Cp�)�|>:���"9N�7�ƈn�v�j�YƷ�@pQy��֑��Q��v!��/K���I�=U�ppDʑ��	V)��:P ��!M��%u�pGG�]1&��ɭ��~1��9��M�}O��$���1Sj����v�� ���0bY�������C 8���(p_X�~'��y߳�l����̕��,,շt:+8.	m��K���[���In��X^v,f�@��8e.���C���Lr��)����2��~���E��<�h�(J)Z�oY��:�x�����ON�jSh^31)�&|s�  mx��iG�N�����C�A�j�3z'��;�+�Ճ�)[��,��T�i55��6q&��7�H�����(0m�E"b��\�B��|r��d,^=ͼ9r=W�_S�\��f��L'{|��d֢=�*G
^�&@4\�}4�o.�#$�W3�$۰~���n�֝��[�.��� U�U�Ŀk!mT,�Vw�����!kL�P�2r *�znX��0�j�uR-����$�9r*Sqa�@Ң.$��N�r��M0.GZ��PVM��
��J�E#x��Kp#7s0sàLF�[B*�!-���Y���ė�j��Y6�]���ľW��D�l�+������fw/\��<�>�{hKR)���8z`�a��O�Jr�t�L>P0N�����/�$�.�?�8�L�͙��zN��q��MI��K��J��njq:���[v'����'�t5�(0
#J�H�}�4�ݜ_�kY�Y�9��n�a��N�N�!�e$�/���]\[�6gq�J�4��w�,Ȍ����kG�ߌ�(��|�����v5 �,kO���'&�s\��5�#�$�냔߆,���ީ7#D��H�{Ě��~��X2��n!�ׁWi�<F/)v~Ģ�v�l��*�$Th�P(�Ѭ�0�-:љ��̨*ܺү�RnkbP>P�?*)ʲ����J�u<P��=����2;�1� �>e]n�R�:����)�	�H*�\r��.�|(gp��L��Y���  ���K�s��������I�M�'G���|��ӄ�����s�!�3�e�3�Bb�H J׮�C�=��5�y��/��w��hWz����J>��{.�;�T7m3Y�x��wo�i|L'sF����V�G�ͤ"'�O��� ��Ž�4��P\��幜��b�R5�����<�*R*�	[Y=	�n�:���$o
��H\�~��'Ō���P��
j-3�����`6,y/|�E�t�����-ia��,o����e�Y��ԈR�	�r0��v���A-ҹw�(<�շe
�(�x�2"t�z:!��c]�j�Z�/64��_15�U������$T�/ճU ��o�QV��Q���d>腲��"ը���l�ӕ��^�����A�~�0�,Z��Ӏ=0���`��ǟ�=����:(�f�H�f���_�+(Q�dK�/�?1K�(@ʌ�?}c�ŀ�j�e���>�Ha�n�����6�(����۷�����"�$R����=<X�
c�8����[��N��<�E��x2�����>����CQ������ʭm���36S(я�A#��ls<����ȊU�'��s�3.D���h~���a���6<
A5:�]V9�J3*j)?� ��!=���>�S>��q2�q�j#\HJ$�z��u���]#\,^��}��*|9H@���EU�V[k�I���g6�[�/
��%n!��$�h�ِ&Yn�34'�����b�9�ƾ��&�#02�-���:���/��2�R|6�ȧ"��GO�C9 �M�&3�A>/��h�Q�!aS��(��F��R!a��=�^�>]��r
)��b�*�pc�~�%E�8Z>`�ZO�j>5���N��I���PH�c|�����ġ��������^�&��3}�����@7����Qo�+��;�.D	T��)�?�P�
��)R�׏!�����eR���aq��%rrg?s��A2���0V��F0zU������w���0��v��=�8ӡ�u��J��g�UJ��"�E<�L�%S�%h��Kɒ�b��nj����"����m z#����t'v��	�7�y�LJ���+�:[1������U9P����2�N%d��d��Y�	#� �5��Z��1���^�"�aD��P���� #v�o�A=_��F�1`x��/��l�ɿ��!��s!ѵ����:Pv_k�`�h�秬�����}Og��{Gy�iKK���`�7+g:��p�泒�f�#�+_v���1J�:i���r,PW~�FA��D�9�)2���m�7��]��U^s�-)I�0����:G�4�b�������"�/_�F�ffՙ��Mu ���!1�_�#�f漻��_��#�����A�ؙ܀�0�����'̴
��'�O1�*u�&�K����.��q����, .Ve�^�|Mx�H�6�4ȸo��k}�����JX���7���<R���$8����E�mp���}�cK�ų�����P�`ܤ�n~!*#�����Ӓ��5G1�Z�<mv�
P���_�c9��вC���Z��L	���'�S��t�!<�V�����iw���p��.!�s�h�;�mbG>9Lf�o���8��?Y<A�

�����KqHn_qܕC�;.C�_�y���>�Ir<L_s��@�@~��#���g�B�ՙD�m���	B���I�=��|��O�L%�EԹlB]%�ɉW�2��M� �.��D!#�w�}�vCK�������x��M�4�;7Lх�=�B���|<J��5m��	ih�wl�(_�>�WpBΈD�������U��3ǙP[k,�f�tn�t|� ���F� ���$De��" �P`>����b�i�Io.�^0ϸ��;��¸�fz�z�^���9j�-�&���G�I����ߗf�� �&|>�3'V�a`Z�?�~�+����o��S�2@���nH���]���
CT���Zs��1D$����!\G�f�Z�\��I�7���{��C_ХB�'��=��!^M�{�=��˗:��es$������	�����?�M��O|�ՍM�!;ʊr:��	Q[����{���h:O�KL'4�G�{ƴΝCŷA�Ge�1�b���}��rwk���{�Fp�zY������J_�+����������~/���'
6�~����/|̈�7F�tqWv�g�F�t ���FGNث��2Aꖚǫ�o���(�J�lJ����\N��H:L�i��@VR�P��K��� �U����1��T��>��T�$b������?������l����9@!��y"@d�m����\�[ЏUq�u� �-/T)5{�8G���~�K�/�YY��7X�D �P,�}������<���'Ղl5�����`%O��J���VO%���*�m��6��N����j%o�$�CE���������r ;�d(�M��cXѾ�1%d���Be-��Z&|��r�P�����d^�)�s�8�ˑɯ;J\f��uКB=R�r� u��ܲ��C��{�����܂2�D������\@ߛh�I��(�M�u��-`g��ݯ�^�	��#�E��$\�$E3l7jLu���47�O@�"����b+kDiG
+$��"�r�ՊI�F-6ڋQFZ.��u"��.5j�[�W�t[�ۋ�-��o���s���������Z�(�PL!�0�������R�um�5X����덦��.C�������Wx�Ś��Շ��m�\3�?�+�hKS�H�d��FmD�j�_O���6�
�,F����[�z���'��F�݃��B��kQ.���� ���t��?x��э��@��g��	��*�ԄX�mͱQTPu9���+Cx��29R$,�K.�){5�.7 �|�2���ܼ�h�<�ܥvJ�i�*& <��!�]b����# �,��<��c=�+k�-C��H�Ϧ�+n�s��g�}���/cV��E��3�������˕ԓ��$��ja�H���$W@B��`�-��TQb��ҜP�PC�1ۂf�I�7�.�))�S(��ϫV��޶�"��*uBHi��W��'�U�}����^Q�Ƽ�6���ƴ�<b���q.�9ca�'B!�������ݏ��m�آI�Z��1�B73xI���I�mt���e�>n၇p��ocJ�%T;
7