��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.f(v����Ih�$,����d�H��zJ���kN-�BA'm��z�:���ϼ��<r`���#���c�,���+b��FO���F����)�f����X8O��Ob�i���Nx�N����;@+�n��O���^u4�'����VP�_m�W,���#D3 ��𕺸�]*�C<�'��LCA]4����]7X:Q���zTԻI^c�����d����VS�����YU� ��)'U�qʱ��H�����h��ŁR{��e��D}�z�_e�b<=ܨ��k�#���'�8W�k@����^� �n�/������,w�2���h�`�$��>�ȼr���+�7���\
��} ���1�^Y@^��Σ���x����f+�_S�Q��Rlp'p��f�c���ʒeˣ��Lv���O��X�n��V��ڛ�,�-�d��QU��@s[Q������M�����|d�;O�"�����<O۔@�l�7��d����Ǉ|u(��roN;�%�PS�BPD���F诋��b�=��O�Q��v4�G�~
��&x�';o��37�?3��S
��y�}�"J*�=˓Y�7?y��Wl��<�;�� ��*̊�����i��������H��1EWX(�k�b1�����ְ-��]�8��7�?��{Ù�pIz+F�H�������_?��6%��p�z,j˧����[���k�M��?ɵF�0ٕo�AZ�z�ܝ�LQ���s��(>ƙ�E�E(�>���ɣ$2���o���WT w!x&d7a�a�Y#) ��xJ��RT`�ld���<�������b�D�-�aͻ!՜Ȥ�Մ�KE�ϝ�q�2��T$L+��K�z��H,�Y8��9�:����t`�_�r�n(HO��v ��(S;�R�~���nqX
����H��n�
ߜ<N��+���9)�Y�Qc������P�`h�2�����>�!~� �>Ek;)�&�RO��9xe�\�����+µ�ϲr���E~u+	ƭ},ok��K 7w��#=� ̶z	X���bp�6���T)GUB%�;��j�}TޓN�L�l:Q�י�f�B�듴�h�۠C������E�,��;�����\ X��졫<l�|lZ��22L��k_	�dX���{�`�w�fL�J���#�жf�r��H��h���]�$a�}a�27@|*b�:����	5_�K�f>�Nt~� ����
U\mWMK*�η�c����Nl4�����!�I��R�+e��ӛ����^q����!�7Bt�Нa(����7n�?�L��ZG�>Ӝ��`2S�C�\MF1�=K>*�ePxT�~@Ǚ��I�6%��x�ѹ8E�W���?����+�9m�N��P赫?�PP��$�jJC�t�'����8�[%�ص	�Pȃ�-u�iyǺh�qd��P��aŗWfǾr�s��� =�t�ܤ��Om�X8بO�p��F�*��e7��!hOoV�I�v���ט�ŋ:�SaMI���g�;��� ��t"}�sb��]���_ G�����ʚ�l��5��P73����?lEgnq�I��,�"���;c6��D�Qϻ�>7TOװxe=qj
�����?�}<ّ��|�;��{n���m�	q��Qm}��G�!O���d���Ǿ�$��4w;��	�W�K���FL��oL�Ed���3Tr,R�����;�����K�jSXq�_�����Y��춡�Ye��������s�z���Y2"4�>�����y�O�dṒ1�P_5[�b��S��$�zs��{���^�V(%i�P�|��g,P��U�8+�R/,��&8��v���.y���b��%~��탪@���pI�_�4�nwv���pLP3�/�Z'�H�j=ٶ�@OWQy��4|�~5/f83>(�61�	�=�����r�c��,��m�+���$w���J�:0&����n.��RG���ۥ��< �y�3D{�q�	��YT4X�׌�oP��c��s��/��^�~��]�ny�L,�Qȥ�ʼ��"�&٩����K*�yC���D�����jQ�{+���&T8���K�|�|�Xʓ#W O_4*+��}�~��/� !
���G�36�AI�Am�ø���E몊\\Y,��Z�g� l�}�0�f�T��E̳��c�,W�~w�s���,��	��M�:��R8w�@oNm�J�46a�a������Kڂ�> �۷4jS����.�lN�F�	�)�ۂ���tٮ�_�_s�$���+g�b�$HUl\*�G��qb�#Ft�jb�̵��eH:�b74��o4��3��>�����B�����+�jD������j=�B@�*�*q&�<�~#pU��hk�s���>΃�_�tN0鿇Lnأ*e���`�B�"���;��`�K�0"=Hq-͌�O)]/mmh�փ�B.ا����r��(ÔuZ?t��:	�DZcxG�){��w/�	�����/2xʑO��J���_��_e����~W��a��٥)|��c���?�?\�g�8��ӡ,��I��xC��e�@���T�t�����u�S��$Jђ���	0q�ۨ����O��M%��Rt�D�SB�Y�� j;��=�,�k	������/�������+��SQ+�o(8���ţ��Z��Am������t��\%]���}zFc�<�0�AS���7[9�6���Ɏ	z!P16m�B�+!g�r���U�j:Z�k#xk Y�۔��揌�=�9[%��+d�k��?�Ήg��Qqc�s��/w]�8��xɅ�B������&�&�=<��]��Mަ�ddٿŞ��= ��é�s��bL:d0�y��g��[�{�v�I�?���>�����W|`�I�E���٣
G-�Fa,y�^Cr�lh�"+�Vy�F��D#����ۛ �CO��$0Mq�3��:!�,���.X�PH�w�KS���(ɖXܛ�"%��N��&�WE5v���+�E���9?;�q8k�/�肌L�B�7)��C2�ʼV�#J	�k{����u�G3@�Q���E��NR��ј�0U���ׂ>F�&0�ѕWm��n��h�x�~ٗZ�h֭]-� /,M��<�Gޠg�9y�S��n�"n O�ae��Q�ǅU�!���w����va�tQ��T�ӝ��&?�Ir{�-ĐR�_��[9�:��������2?�A�:���RІ�&*����?��5L����?��K7\�$�3�=
�n���@���A��y��1��0�������R{�::eLY,�*�_+�a �?���fz�Yi̧j;LD�ϗ�U���'�8��x5	�3�`�8�⭠f���+���2�r��)�<b�k�~����l��ד�Rj}%�bEa^�@P�N���,�ǚ8gqI]�#B����xœQ;X��O��%�W���I��@�<���J: 2ߞ�wih/>�Y$��3��-��.����l��M�BC��J���iI���� ��m��OH�����7���p��e�6��-9=��uT��1�����I�9F��ƍ��#�f��D��j�qٰN����E)b�q!��Ê,g��ӕ�'�caw��0�v�V��6v���a������a�B�]�:��8T�!���<%M�`3�b`L��L>dA�bBG�v��A��f����@;:�q�؜�~����֛F��:�����"}�o��;���X�`P9u��?d�'��㣿�K�,�G��1c(�S*�Kױ&+v��wR�8�q�߹٪{���i�ݑ�� g4{�>�����mw��9�?����lE���>�V���x�����T��O|�.F�j�G^�s9�������K�5T�D�W�g��_0e���3���z`��fZ�� _��~�>���ݑ|6n� �%W��9�'������&X����z���E\�g��"{��K�����(wFFIG��H?�朐� ��d�yeܼ� a��G�����qy.Uȧ#BZ��L��l�ك�$+�qu���@)GXF�{�֧z�=�7r,�M�Z�.-QG<͕�-t�.��"��i�h��^�2�Y��N�e��,s�����Y�L乃D;��(���=e�_)oL�'�+^�wI���Yg�e��<J�q���J��*c�#��������P*g�-��i"˶��6�5>����v(h�D-��,�Ѿw�>����b�w��M=��)n�g��We�o�Y[D>�j-��a���a�tк-���,p*h�T��|)�u������C[�]e�!�'a��nt�qY�G�S���Z�$�\y�R��sҚ�����ŪN;}PB,�EU����T�  ��N7�j��1�_��:�$?u�g3Z�7c�8�9tJZ�I�1�E��>�8�A��퀡��=p��H���?(ix�D�+��[�=u�^V�-F�m��>��6���U��M��"qG̡Naz�E慄6��w,��R��s��x�>::�a�Q90�Z�=���m�d���jrLSh����i� �-q��F���\�O��X�7���D�%����@>=��0��Er�/�����27����O�\բ�:kq�.d�6�_B�[y���/�������Z1x^kT���O#�!�(����^t'���Mu	�Y²S9�CQ�c�#�U�;�� s���5:�)�:l&���ݮ�]�O�����b������缾�D��3�%�Vm�~��=�܀75�w%���'w;_B��$Y�"�S�'�S�u���T�]�t�kN��M̻[���)��I)�	�1:2�G�n�_��sfԔt���L�K����9�a�ss�}�{���'��Ghy�f�ͣ��p|�n�L��x�a�z���P�-\^��fD�T�<�{��qXغ'ڮ��y�Ev :|'o�	적�B36 �����wad�jOQ��4D�Q��{A �E#C�����������s[���{�:�~�#�i5����i���+a�/�d�%Dܨ��k'�C�]���tx�
�X`�Ĵ��+E���/P�أBpՉKU����l[�A'�	%7!ky�����G7�p=�Յ�\đyw�k��^VD-���&D����,�J��2Y���-��E�Èw���K�2c�i7S[9���rPG=�Sǝ�A�!����yLO4��)Z�8�������Ћ�� l�>�jo}h�+|�R	���ʜ�ɭi�@�