��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.f(v����IC�ݟ��OTӌ[H'#���S�z�4��J+@�b����	jȕT��/�¹��#��P#�)���%$:���M�s�Ml��,=�z �OU���#��Gn"}N�s�-���r�3а�-�@��I?�ȕ@\��.�+}j2ON<�&[����o�<��=mҪ�/�`=<���X��7|�����(��c��AYd��D<�����c��ۄQ1�X�V�8���4���,Y����GgI_ؿk���c�^�c�&�WZ� ��)�ܤSFK*�Q�%e�=��{����mi?ҝ���ݢ��}?����嗌�?�_ϋ��� m�n���*<m�5樫)��e	�\
;=t���˂��%����.����߁��b������GxB�b,*�pA3�a]���Q���u����s���$�l�ĕE?�h{oH+$q���P��#09��}��܃;&�Kn�A$�	{-��oy��5ے�[����x�(��h֤r���!<��o���$s��NS9':����|&p�مd�&���":vm�b��&q�׻��4�5���$�H��.8���H�>J�W�� &�'���h�:0Q�e	Inp&G#V�^���q+����R�*;�p����Q��Q�Ƿt޸K��3�a�A��V���f��c�8ɫQ)�Vݓ�n��C\��6�s��72M{%���v^�`�Lw�rJ���%�Ukn"���,���f+V�H��w��Ҝ�W�e+����3P���i��3J�����D佊��F��ղ
e����z��a�[�o�{9loGO��\P����Ҧ���_��=V=j���L������ְCگ�{��[�/]1��+6�/��6����[�#V����P���/�p�̶��}�X�C��G(��T�NT�/�:Uƺ	�:�
n�E�K��j�F��uo�1���V�ηrγ�茵�m���hu0���R�{S�cR�@](5g���$o���7�K�����6�\'��[��	/P��������.:����+~�F��f%�[t�]d��e]6�t�����ۻo Ψ��#�즾�RK��1	��!�_�,hx��;*�C����ݩ��N��+�ݣ����%�r�!<v�p٣~/�b�m��Wi�oBkux��y��8�{r��o9����e�*��|��%އ���Y�k�����;���pBg��o�|� �
��s�р�����߯�'.e�>�J�k�Р8j	�S�����8����5�4��/�ޑ��������T.�8�Y���C�����_槴:� ��t�үmf+����=`��|��t����>�S:}�(��J쉄� ���An��;�,Z�B�
B���ʂ�%�:�����A�;a�?��1��}�.�̠��/���}V:�3�����˥\�]���70;&S�H)e�"&n�@9�+ ��5A�߫xF��*c^znC-���w;ɡ��T�c>��4x��Z�r6�%��t�8,+K�s��������}���N�o;�0w+���D%�^М ى������>�T�4�~2�+H`u����c�=)�W�ɧ�wq}��hSLo���0��&�$)~�k�i�PS͈���;����c����q;��1�Bq{�QI�Eeu�n:��[�����N���.�"��@S1�%k9�e�@U�<�2�.<��O��yG�	mY��u��d��p�#�]>�����^S�<����_��>�X��:�;��$�ö�5'V���Q�=���s�`݊��q;���OJ�n$�&"�jݒ	|�&�D��Ḱ����j�0�����I��}���W�ٖ!�\5`��ʲ\��o�p����3����c&�@�x+Ё��;uσ��;~kJ9}��b%E�ȝ>	c6��@�v)��d��|�"��c��h�R�ϔ��B"E=ߟL��X�!����&Y@濍��B�/g$�o��h�,�#∓(y�~�����&=G���ӧ��?aJ����@���I�����g���1�x^���
	�"//�bX{�3��������I&�^����޺�����gI�2�(��)1�R��o��7K��E&@��#�a��<J��1T���&\�� ��Eԩ:�$��d��=�+X��77ò���9�<�B��,g�&���zNr�gќo��fVC+�`�ac[�7�Y쩆�l���ɐ+7����T�}%��^�t9�vi̊	V�!$_N�k8o`�g��_�1��C֍�{W�E��Ė�ꍷs�a �d�8Ԗ6��To��$Pt�O�XA+�"��Ɩ_7wl�Lx��,Ľ�)s�6�� �{�J.�;�:����B�"�yr)�ά7"9�n��3��XR
P;�*�������.�ӵP�3�K����E���\g�!<P�a�1&���=ب)�s�H� �lc��t����b�Y��~��2��rGf�@1�Ѝ�x�'㑆vݖ�f���s���,Q��u���,�	_��K�mp�0;����ނ�O15g*�h&����T�㋄-ndT3�.��FY�)��&9�>L�t%;4f��+J'cwqSh�w��2F���[�$m�N�L	,$�5TF����I�olC˽NKN9�:�6隞�\�	�wH�v�f`�!�wX;�1����w-xY�?�r��KBÂ�%�S��0V�@zB�!�c{�B,�}���F㻟44Ӯ��@)��jDT�a��/n�ǎ�H1ַ�W��gn�0�+-�x�k�ޕ��q��τ�����S���8�z4�K�6Y�u���0��(P(���h��z����v�uP�X~`/gݥ��7�8d>�͕��ss�LOM˴��e?����ι���C�T��m�RG�
��h���Bg\�np���Yz4��N���Ɐ�o���:YܼHܭ*�6یH����H������FPg��^?Z�gq�Ǥ��÷j�� z��ٮ�;�HH\>T����-����1��o�'\iG	h8�\Տ�~aΈ*SK��o��������{$�vu2[S�RحȺ�I �Y�b�Ds������_��N{KAU
3n;��L�����V.XM��`h�6p�D�>�?W?�
��g�r���b q����V��e�� N`
7���
i��2��1HH����(�Ent�pK+��X�?��G��ÚT��h��ѣ?��[�H���2BN/np��&no�9!rƐ�7�����x]G>�9��F��Op�1D��n�K�oϋ������3`{:�e��ׄC��!��Z�$m尿o�׹C&v��	�7wr.�~� q!t�r����3G�Uc8|�ߍ3�*3V�-ο�o>�F2?�,-��=WH��<~f��U��&���_X�X^A�����.r���6�U���ja_.I����,W:��8[p�(!�@2�� ���hu-�嚖0�F\j��#i���*�L	J�Ғ�Ļ�\�����N����	��gipw�)*v�"6���n��p�G���kH�m�=NH�	;��-�q�&�'�^�HwH���;���g<���.�ѻۡ�A�s����O�L��i.�ѵ��R(���eX���C��]O�qy��2��+v��w���0�t�㓟a�����0�����"����f-2L��\��f��D ����8���O���d7�'+-���G¶�G�T!WH��6R�Q�<|Y@������&N�^4����S�rjP�(���JB�1�E��U���;�sI��`�ĥ��^��a��20�2F�':���<�^�B��]��sv,���q\)�7�Ĥ�`q�:�p�� �����ķ�6ښw/@S�l8�[ϻpx�k�SN����8�H�'6ztf�@�j]D�K���#@>��r��R]HڇP}c᳽�r��r��G�WK̓58�"��0��w��S��6�,>�?�m)}�V7V���#=����G�1���።�`Nz�c��,�Gl�w]����=�i�*Pv��H�	��V�0G���>[����)_�"J�x��/4�
��N�|�U��K��T2�<�C�'ߞ!
���b��/r�A#C��ǽW{�1+����zb��ǪL5�R
Q&y�0�M�~�/��LNoj�C,9hA7�RI$�m�<�?#�f�̓+Q��[ϊ���~����{TK��+#����;�Cy^�V�_yp˴���VI�i�>�ֆp�ė2�3e�{Ŷ��F��\s�W��Q�%~CT�ɑ��q��J3��|��h�Cm
� �3q.��K3�	ěe�a�T��E?���U�(������V�n}CE-��7��-�b8/�S�Q�`5o����ւз	��K�t�`����`����W�s����w��\�<&$��I�ΨjP���Q&J�u�CypF8(p�ڵ�S���J� �?����N�6��"	����Їx�K�X�B�����e��Uf�� R��:Nb��0�d_�b�W��-��WK��9��*$��[Nt��$�[�0���oE���u>x�a ��G�qZ�����V�D�F�k��i�3]:����2��?���/�c*)Hw��w�'���V�1���p5h��\�7:����tb]s�#�W�"�D{|�jF<H����#V`n̝d�ΌfP8H�$@�|g8��;O>�*�n��q�5Yr�h�S�ӫ�HD��F�\��o^j�z�H�I�NF��_��]]�q�����c&^\��0�LK�)�oi{�k�Wz	mO��V�Ja����7�k������4f.�=�V���F�QsHlF��6�Ĩ��d��NΛ�'�"?�-I�nIc�8襢H�����V#g��ZHFH���,Fga}u6L�ä�FaY��UD��"M��Y���e� �6`�� �l�G-�yة�[U)w]~�ʿzI����54#�)i�F�tNHY��2'V�q�� @� .u��3c�M >�Nj�QJ������Q�ip�q����QW�Gt	˹�Z�����L�����@:��D�_9�?|���HhMQ��}c����s��ث�?aN�Ҟ�P��xRܙXm7\'~�,W +
���^*��P�`�゚ͩ(�n�h�ܕ*��= '�x��x^JT"ʭ̓��|K�I�
mh���.��[�%v���Q�g\�5�Z4{�=���b2A�-�㥓����iw�俇�8��XY�G(���D�0m�iP�e��[�[S.�f!=�tJ\	�ezۄ�"$G_`M{���Y���ՑXR�Zit�9�|��w�D�S,p�չY�}8�K��}LV�0�v�_9Ĉ�?j���œ���g\��}��o�s! A�f�ql�,�Q$�>��ج��&�Ы�sљB9�4%T�M$|�����u1�b+7�(B"o��xV� ��=޻6�Os�+� ��rt׏1� K�6�lH����S�߾O��rv�T �<1|�Q5s}���A��_�
L	ZP�ek��K��'��}���j�^�$�ATL��_`��At���3?) �휹�b0"YB�Ԝ�\\1V	��赀 �&�L���O��\G���������N�P�N��^� i8ui�$pl��`�E���-��<��
z�y���~;0��py��_����C��qZ_��m&d	�mÃԸM_T�2e�V��n>X�"_����V+�f/%��